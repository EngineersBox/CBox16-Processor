//  A testbench for control_unit_RS2_tb
`timescale 1us/1ns

module control_unit_RS2_tb;
    reg [15:0] INST;
    wire [1:0] ALUOP;
    wire [2:0] RS1;
    wire [2:0] RS2;
    wire [2:0] WS;
    wire STR;
    wire WE;
    wire [1:0] DMUX;
    wire LDR;

  control_unit control_unit0 (
    .INST(INST),
    .ALUOP(ALUOP),
    .RS1(RS1),
    .RS2(RS2),
    .WS(WS),
    .STR(STR),
    .WE(WE),
    .DMUX(DMUX),
    .LDR(LDR)
  );

    reg [18:0] patterns[0:2559];
    integer i;

    initial begin
      patterns[0] = 19'b1000000000000000_000;
      patterns[1] = 19'b1001000000000000_000;
      patterns[2] = 19'b1010000000000000_000;
      patterns[3] = 19'b1011000000000000_000;
      patterns[4] = 19'b0100000000000000_000;
      patterns[5] = 19'b1000000000000001_001;
      patterns[6] = 19'b1001000000000001_001;
      patterns[7] = 19'b1010000000000001_001;
      patterns[8] = 19'b1011000000000001_001;
      patterns[9] = 19'b0100000000000000_000;
      patterns[10] = 19'b1000000000000010_010;
      patterns[11] = 19'b1001000000000010_010;
      patterns[12] = 19'b1010000000000010_010;
      patterns[13] = 19'b1011000000000010_010;
      patterns[14] = 19'b0100000000000000_000;
      patterns[15] = 19'b1000000000000011_011;
      patterns[16] = 19'b1001000000000011_011;
      patterns[17] = 19'b1010000000000011_011;
      patterns[18] = 19'b1011000000000011_011;
      patterns[19] = 19'b0100000000000000_000;
      patterns[20] = 19'b1000000000000100_100;
      patterns[21] = 19'b1001000000000100_100;
      patterns[22] = 19'b1010000000000100_100;
      patterns[23] = 19'b1011000000000100_100;
      patterns[24] = 19'b0100000000000000_000;
      patterns[25] = 19'b1000000000000101_101;
      patterns[26] = 19'b1001000000000101_101;
      patterns[27] = 19'b1010000000000101_101;
      patterns[28] = 19'b1011000000000101_101;
      patterns[29] = 19'b0100000000000000_000;
      patterns[30] = 19'b1000000000000110_110;
      patterns[31] = 19'b1001000000000110_110;
      patterns[32] = 19'b1010000000000110_110;
      patterns[33] = 19'b1011000000000110_110;
      patterns[34] = 19'b0100000000000000_000;
      patterns[35] = 19'b1000000000000111_111;
      patterns[36] = 19'b1001000000000111_111;
      patterns[37] = 19'b1010000000000111_111;
      patterns[38] = 19'b1011000000000111_111;
      patterns[39] = 19'b0100000000000000_000;
      patterns[40] = 19'b1000000000010000_000;
      patterns[41] = 19'b1001000000010000_000;
      patterns[42] = 19'b1010000000010000_000;
      patterns[43] = 19'b1011000000010000_000;
      patterns[44] = 19'b0100000000010000_000;
      patterns[45] = 19'b1000000000010001_001;
      patterns[46] = 19'b1001000000010001_001;
      patterns[47] = 19'b1010000000010001_001;
      patterns[48] = 19'b1011000000010001_001;
      patterns[49] = 19'b0100000000010000_000;
      patterns[50] = 19'b1000000000010010_010;
      patterns[51] = 19'b1001000000010010_010;
      patterns[52] = 19'b1010000000010010_010;
      patterns[53] = 19'b1011000000010010_010;
      patterns[54] = 19'b0100000000010000_000;
      patterns[55] = 19'b1000000000010011_011;
      patterns[56] = 19'b1001000000010011_011;
      patterns[57] = 19'b1010000000010011_011;
      patterns[58] = 19'b1011000000010011_011;
      patterns[59] = 19'b0100000000010000_000;
      patterns[60] = 19'b1000000000010100_100;
      patterns[61] = 19'b1001000000010100_100;
      patterns[62] = 19'b1010000000010100_100;
      patterns[63] = 19'b1011000000010100_100;
      patterns[64] = 19'b0100000000010000_000;
      patterns[65] = 19'b1000000000010101_101;
      patterns[66] = 19'b1001000000010101_101;
      patterns[67] = 19'b1010000000010101_101;
      patterns[68] = 19'b1011000000010101_101;
      patterns[69] = 19'b0100000000010000_000;
      patterns[70] = 19'b1000000000010110_110;
      patterns[71] = 19'b1001000000010110_110;
      patterns[72] = 19'b1010000000010110_110;
      patterns[73] = 19'b1011000000010110_110;
      patterns[74] = 19'b0100000000010000_000;
      patterns[75] = 19'b1000000000010111_111;
      patterns[76] = 19'b1001000000010111_111;
      patterns[77] = 19'b1010000000010111_111;
      patterns[78] = 19'b1011000000010111_111;
      patterns[79] = 19'b0100000000010000_000;
      patterns[80] = 19'b1000000000100000_000;
      patterns[81] = 19'b1001000000100000_000;
      patterns[82] = 19'b1010000000100000_000;
      patterns[83] = 19'b1011000000100000_000;
      patterns[84] = 19'b0100000000100000_000;
      patterns[85] = 19'b1000000000100001_001;
      patterns[86] = 19'b1001000000100001_001;
      patterns[87] = 19'b1010000000100001_001;
      patterns[88] = 19'b1011000000100001_001;
      patterns[89] = 19'b0100000000100000_000;
      patterns[90] = 19'b1000000000100010_010;
      patterns[91] = 19'b1001000000100010_010;
      patterns[92] = 19'b1010000000100010_010;
      patterns[93] = 19'b1011000000100010_010;
      patterns[94] = 19'b0100000000100000_000;
      patterns[95] = 19'b1000000000100011_011;
      patterns[96] = 19'b1001000000100011_011;
      patterns[97] = 19'b1010000000100011_011;
      patterns[98] = 19'b1011000000100011_011;
      patterns[99] = 19'b0100000000100000_000;
      patterns[100] = 19'b1000000000100100_100;
      patterns[101] = 19'b1001000000100100_100;
      patterns[102] = 19'b1010000000100100_100;
      patterns[103] = 19'b1011000000100100_100;
      patterns[104] = 19'b0100000000100000_000;
      patterns[105] = 19'b1000000000100101_101;
      patterns[106] = 19'b1001000000100101_101;
      patterns[107] = 19'b1010000000100101_101;
      patterns[108] = 19'b1011000000100101_101;
      patterns[109] = 19'b0100000000100000_000;
      patterns[110] = 19'b1000000000100110_110;
      patterns[111] = 19'b1001000000100110_110;
      patterns[112] = 19'b1010000000100110_110;
      patterns[113] = 19'b1011000000100110_110;
      patterns[114] = 19'b0100000000100000_000;
      patterns[115] = 19'b1000000000100111_111;
      patterns[116] = 19'b1001000000100111_111;
      patterns[117] = 19'b1010000000100111_111;
      patterns[118] = 19'b1011000000100111_111;
      patterns[119] = 19'b0100000000100000_000;
      patterns[120] = 19'b1000000000110000_000;
      patterns[121] = 19'b1001000000110000_000;
      patterns[122] = 19'b1010000000110000_000;
      patterns[123] = 19'b1011000000110000_000;
      patterns[124] = 19'b0100000000110000_000;
      patterns[125] = 19'b1000000000110001_001;
      patterns[126] = 19'b1001000000110001_001;
      patterns[127] = 19'b1010000000110001_001;
      patterns[128] = 19'b1011000000110001_001;
      patterns[129] = 19'b0100000000110000_000;
      patterns[130] = 19'b1000000000110010_010;
      patterns[131] = 19'b1001000000110010_010;
      patterns[132] = 19'b1010000000110010_010;
      patterns[133] = 19'b1011000000110010_010;
      patterns[134] = 19'b0100000000110000_000;
      patterns[135] = 19'b1000000000110011_011;
      patterns[136] = 19'b1001000000110011_011;
      patterns[137] = 19'b1010000000110011_011;
      patterns[138] = 19'b1011000000110011_011;
      patterns[139] = 19'b0100000000110000_000;
      patterns[140] = 19'b1000000000110100_100;
      patterns[141] = 19'b1001000000110100_100;
      patterns[142] = 19'b1010000000110100_100;
      patterns[143] = 19'b1011000000110100_100;
      patterns[144] = 19'b0100000000110000_000;
      patterns[145] = 19'b1000000000110101_101;
      patterns[146] = 19'b1001000000110101_101;
      patterns[147] = 19'b1010000000110101_101;
      patterns[148] = 19'b1011000000110101_101;
      patterns[149] = 19'b0100000000110000_000;
      patterns[150] = 19'b1000000000110110_110;
      patterns[151] = 19'b1001000000110110_110;
      patterns[152] = 19'b1010000000110110_110;
      patterns[153] = 19'b1011000000110110_110;
      patterns[154] = 19'b0100000000110000_000;
      patterns[155] = 19'b1000000000110111_111;
      patterns[156] = 19'b1001000000110111_111;
      patterns[157] = 19'b1010000000110111_111;
      patterns[158] = 19'b1011000000110111_111;
      patterns[159] = 19'b0100000000110000_000;
      patterns[160] = 19'b1000000001000000_000;
      patterns[161] = 19'b1001000001000000_000;
      patterns[162] = 19'b1010000001000000_000;
      patterns[163] = 19'b1011000001000000_000;
      patterns[164] = 19'b0100000001000000_000;
      patterns[165] = 19'b1000000001000001_001;
      patterns[166] = 19'b1001000001000001_001;
      patterns[167] = 19'b1010000001000001_001;
      patterns[168] = 19'b1011000001000001_001;
      patterns[169] = 19'b0100000001000000_000;
      patterns[170] = 19'b1000000001000010_010;
      patterns[171] = 19'b1001000001000010_010;
      patterns[172] = 19'b1010000001000010_010;
      patterns[173] = 19'b1011000001000010_010;
      patterns[174] = 19'b0100000001000000_000;
      patterns[175] = 19'b1000000001000011_011;
      patterns[176] = 19'b1001000001000011_011;
      patterns[177] = 19'b1010000001000011_011;
      patterns[178] = 19'b1011000001000011_011;
      patterns[179] = 19'b0100000001000000_000;
      patterns[180] = 19'b1000000001000100_100;
      patterns[181] = 19'b1001000001000100_100;
      patterns[182] = 19'b1010000001000100_100;
      patterns[183] = 19'b1011000001000100_100;
      patterns[184] = 19'b0100000001000000_000;
      patterns[185] = 19'b1000000001000101_101;
      patterns[186] = 19'b1001000001000101_101;
      patterns[187] = 19'b1010000001000101_101;
      patterns[188] = 19'b1011000001000101_101;
      patterns[189] = 19'b0100000001000000_000;
      patterns[190] = 19'b1000000001000110_110;
      patterns[191] = 19'b1001000001000110_110;
      patterns[192] = 19'b1010000001000110_110;
      patterns[193] = 19'b1011000001000110_110;
      patterns[194] = 19'b0100000001000000_000;
      patterns[195] = 19'b1000000001000111_111;
      patterns[196] = 19'b1001000001000111_111;
      patterns[197] = 19'b1010000001000111_111;
      patterns[198] = 19'b1011000001000111_111;
      patterns[199] = 19'b0100000001000000_000;
      patterns[200] = 19'b1000000001010000_000;
      patterns[201] = 19'b1001000001010000_000;
      patterns[202] = 19'b1010000001010000_000;
      patterns[203] = 19'b1011000001010000_000;
      patterns[204] = 19'b0100000001010000_000;
      patterns[205] = 19'b1000000001010001_001;
      patterns[206] = 19'b1001000001010001_001;
      patterns[207] = 19'b1010000001010001_001;
      patterns[208] = 19'b1011000001010001_001;
      patterns[209] = 19'b0100000001010000_000;
      patterns[210] = 19'b1000000001010010_010;
      patterns[211] = 19'b1001000001010010_010;
      patterns[212] = 19'b1010000001010010_010;
      patterns[213] = 19'b1011000001010010_010;
      patterns[214] = 19'b0100000001010000_000;
      patterns[215] = 19'b1000000001010011_011;
      patterns[216] = 19'b1001000001010011_011;
      patterns[217] = 19'b1010000001010011_011;
      patterns[218] = 19'b1011000001010011_011;
      patterns[219] = 19'b0100000001010000_000;
      patterns[220] = 19'b1000000001010100_100;
      patterns[221] = 19'b1001000001010100_100;
      patterns[222] = 19'b1010000001010100_100;
      patterns[223] = 19'b1011000001010100_100;
      patterns[224] = 19'b0100000001010000_000;
      patterns[225] = 19'b1000000001010101_101;
      patterns[226] = 19'b1001000001010101_101;
      patterns[227] = 19'b1010000001010101_101;
      patterns[228] = 19'b1011000001010101_101;
      patterns[229] = 19'b0100000001010000_000;
      patterns[230] = 19'b1000000001010110_110;
      patterns[231] = 19'b1001000001010110_110;
      patterns[232] = 19'b1010000001010110_110;
      patterns[233] = 19'b1011000001010110_110;
      patterns[234] = 19'b0100000001010000_000;
      patterns[235] = 19'b1000000001010111_111;
      patterns[236] = 19'b1001000001010111_111;
      patterns[237] = 19'b1010000001010111_111;
      patterns[238] = 19'b1011000001010111_111;
      patterns[239] = 19'b0100000001010000_000;
      patterns[240] = 19'b1000000001100000_000;
      patterns[241] = 19'b1001000001100000_000;
      patterns[242] = 19'b1010000001100000_000;
      patterns[243] = 19'b1011000001100000_000;
      patterns[244] = 19'b0100000001100000_000;
      patterns[245] = 19'b1000000001100001_001;
      patterns[246] = 19'b1001000001100001_001;
      patterns[247] = 19'b1010000001100001_001;
      patterns[248] = 19'b1011000001100001_001;
      patterns[249] = 19'b0100000001100000_000;
      patterns[250] = 19'b1000000001100010_010;
      patterns[251] = 19'b1001000001100010_010;
      patterns[252] = 19'b1010000001100010_010;
      patterns[253] = 19'b1011000001100010_010;
      patterns[254] = 19'b0100000001100000_000;
      patterns[255] = 19'b1000000001100011_011;
      patterns[256] = 19'b1001000001100011_011;
      patterns[257] = 19'b1010000001100011_011;
      patterns[258] = 19'b1011000001100011_011;
      patterns[259] = 19'b0100000001100000_000;
      patterns[260] = 19'b1000000001100100_100;
      patterns[261] = 19'b1001000001100100_100;
      patterns[262] = 19'b1010000001100100_100;
      patterns[263] = 19'b1011000001100100_100;
      patterns[264] = 19'b0100000001100000_000;
      patterns[265] = 19'b1000000001100101_101;
      patterns[266] = 19'b1001000001100101_101;
      patterns[267] = 19'b1010000001100101_101;
      patterns[268] = 19'b1011000001100101_101;
      patterns[269] = 19'b0100000001100000_000;
      patterns[270] = 19'b1000000001100110_110;
      patterns[271] = 19'b1001000001100110_110;
      patterns[272] = 19'b1010000001100110_110;
      patterns[273] = 19'b1011000001100110_110;
      patterns[274] = 19'b0100000001100000_000;
      patterns[275] = 19'b1000000001100111_111;
      patterns[276] = 19'b1001000001100111_111;
      patterns[277] = 19'b1010000001100111_111;
      patterns[278] = 19'b1011000001100111_111;
      patterns[279] = 19'b0100000001100000_000;
      patterns[280] = 19'b1000000001110000_000;
      patterns[281] = 19'b1001000001110000_000;
      patterns[282] = 19'b1010000001110000_000;
      patterns[283] = 19'b1011000001110000_000;
      patterns[284] = 19'b0100000001110000_000;
      patterns[285] = 19'b1000000001110001_001;
      patterns[286] = 19'b1001000001110001_001;
      patterns[287] = 19'b1010000001110001_001;
      patterns[288] = 19'b1011000001110001_001;
      patterns[289] = 19'b0100000001110000_000;
      patterns[290] = 19'b1000000001110010_010;
      patterns[291] = 19'b1001000001110010_010;
      patterns[292] = 19'b1010000001110010_010;
      patterns[293] = 19'b1011000001110010_010;
      patterns[294] = 19'b0100000001110000_000;
      patterns[295] = 19'b1000000001110011_011;
      patterns[296] = 19'b1001000001110011_011;
      patterns[297] = 19'b1010000001110011_011;
      patterns[298] = 19'b1011000001110011_011;
      patterns[299] = 19'b0100000001110000_000;
      patterns[300] = 19'b1000000001110100_100;
      patterns[301] = 19'b1001000001110100_100;
      patterns[302] = 19'b1010000001110100_100;
      patterns[303] = 19'b1011000001110100_100;
      patterns[304] = 19'b0100000001110000_000;
      patterns[305] = 19'b1000000001110101_101;
      patterns[306] = 19'b1001000001110101_101;
      patterns[307] = 19'b1010000001110101_101;
      patterns[308] = 19'b1011000001110101_101;
      patterns[309] = 19'b0100000001110000_000;
      patterns[310] = 19'b1000000001110110_110;
      patterns[311] = 19'b1001000001110110_110;
      patterns[312] = 19'b1010000001110110_110;
      patterns[313] = 19'b1011000001110110_110;
      patterns[314] = 19'b0100000001110000_000;
      patterns[315] = 19'b1000000001110111_111;
      patterns[316] = 19'b1001000001110111_111;
      patterns[317] = 19'b1010000001110111_111;
      patterns[318] = 19'b1011000001110111_111;
      patterns[319] = 19'b0100000001110000_000;
      patterns[320] = 19'b1000000100000000_000;
      patterns[321] = 19'b1001000100000000_000;
      patterns[322] = 19'b1010000100000000_000;
      patterns[323] = 19'b1011000100000000_000;
      patterns[324] = 19'b0100000100000000_001;
      patterns[325] = 19'b1000000100000001_001;
      patterns[326] = 19'b1001000100000001_001;
      patterns[327] = 19'b1010000100000001_001;
      patterns[328] = 19'b1011000100000001_001;
      patterns[329] = 19'b0100000100000000_001;
      patterns[330] = 19'b1000000100000010_010;
      patterns[331] = 19'b1001000100000010_010;
      patterns[332] = 19'b1010000100000010_010;
      patterns[333] = 19'b1011000100000010_010;
      patterns[334] = 19'b0100000100000000_001;
      patterns[335] = 19'b1000000100000011_011;
      patterns[336] = 19'b1001000100000011_011;
      patterns[337] = 19'b1010000100000011_011;
      patterns[338] = 19'b1011000100000011_011;
      patterns[339] = 19'b0100000100000000_001;
      patterns[340] = 19'b1000000100000100_100;
      patterns[341] = 19'b1001000100000100_100;
      patterns[342] = 19'b1010000100000100_100;
      patterns[343] = 19'b1011000100000100_100;
      patterns[344] = 19'b0100000100000000_001;
      patterns[345] = 19'b1000000100000101_101;
      patterns[346] = 19'b1001000100000101_101;
      patterns[347] = 19'b1010000100000101_101;
      patterns[348] = 19'b1011000100000101_101;
      patterns[349] = 19'b0100000100000000_001;
      patterns[350] = 19'b1000000100000110_110;
      patterns[351] = 19'b1001000100000110_110;
      patterns[352] = 19'b1010000100000110_110;
      patterns[353] = 19'b1011000100000110_110;
      patterns[354] = 19'b0100000100000000_001;
      patterns[355] = 19'b1000000100000111_111;
      patterns[356] = 19'b1001000100000111_111;
      patterns[357] = 19'b1010000100000111_111;
      patterns[358] = 19'b1011000100000111_111;
      patterns[359] = 19'b0100000100000000_001;
      patterns[360] = 19'b1000000100010000_000;
      patterns[361] = 19'b1001000100010000_000;
      patterns[362] = 19'b1010000100010000_000;
      patterns[363] = 19'b1011000100010000_000;
      patterns[364] = 19'b0100000100010000_001;
      patterns[365] = 19'b1000000100010001_001;
      patterns[366] = 19'b1001000100010001_001;
      patterns[367] = 19'b1010000100010001_001;
      patterns[368] = 19'b1011000100010001_001;
      patterns[369] = 19'b0100000100010000_001;
      patterns[370] = 19'b1000000100010010_010;
      patterns[371] = 19'b1001000100010010_010;
      patterns[372] = 19'b1010000100010010_010;
      patterns[373] = 19'b1011000100010010_010;
      patterns[374] = 19'b0100000100010000_001;
      patterns[375] = 19'b1000000100010011_011;
      patterns[376] = 19'b1001000100010011_011;
      patterns[377] = 19'b1010000100010011_011;
      patterns[378] = 19'b1011000100010011_011;
      patterns[379] = 19'b0100000100010000_001;
      patterns[380] = 19'b1000000100010100_100;
      patterns[381] = 19'b1001000100010100_100;
      patterns[382] = 19'b1010000100010100_100;
      patterns[383] = 19'b1011000100010100_100;
      patterns[384] = 19'b0100000100010000_001;
      patterns[385] = 19'b1000000100010101_101;
      patterns[386] = 19'b1001000100010101_101;
      patterns[387] = 19'b1010000100010101_101;
      patterns[388] = 19'b1011000100010101_101;
      patterns[389] = 19'b0100000100010000_001;
      patterns[390] = 19'b1000000100010110_110;
      patterns[391] = 19'b1001000100010110_110;
      patterns[392] = 19'b1010000100010110_110;
      patterns[393] = 19'b1011000100010110_110;
      patterns[394] = 19'b0100000100010000_001;
      patterns[395] = 19'b1000000100010111_111;
      patterns[396] = 19'b1001000100010111_111;
      patterns[397] = 19'b1010000100010111_111;
      patterns[398] = 19'b1011000100010111_111;
      patterns[399] = 19'b0100000100010000_001;
      patterns[400] = 19'b1000000100100000_000;
      patterns[401] = 19'b1001000100100000_000;
      patterns[402] = 19'b1010000100100000_000;
      patterns[403] = 19'b1011000100100000_000;
      patterns[404] = 19'b0100000100100000_001;
      patterns[405] = 19'b1000000100100001_001;
      patterns[406] = 19'b1001000100100001_001;
      patterns[407] = 19'b1010000100100001_001;
      patterns[408] = 19'b1011000100100001_001;
      patterns[409] = 19'b0100000100100000_001;
      patterns[410] = 19'b1000000100100010_010;
      patterns[411] = 19'b1001000100100010_010;
      patterns[412] = 19'b1010000100100010_010;
      patterns[413] = 19'b1011000100100010_010;
      patterns[414] = 19'b0100000100100000_001;
      patterns[415] = 19'b1000000100100011_011;
      patterns[416] = 19'b1001000100100011_011;
      patterns[417] = 19'b1010000100100011_011;
      patterns[418] = 19'b1011000100100011_011;
      patterns[419] = 19'b0100000100100000_001;
      patterns[420] = 19'b1000000100100100_100;
      patterns[421] = 19'b1001000100100100_100;
      patterns[422] = 19'b1010000100100100_100;
      patterns[423] = 19'b1011000100100100_100;
      patterns[424] = 19'b0100000100100000_001;
      patterns[425] = 19'b1000000100100101_101;
      patterns[426] = 19'b1001000100100101_101;
      patterns[427] = 19'b1010000100100101_101;
      patterns[428] = 19'b1011000100100101_101;
      patterns[429] = 19'b0100000100100000_001;
      patterns[430] = 19'b1000000100100110_110;
      patterns[431] = 19'b1001000100100110_110;
      patterns[432] = 19'b1010000100100110_110;
      patterns[433] = 19'b1011000100100110_110;
      patterns[434] = 19'b0100000100100000_001;
      patterns[435] = 19'b1000000100100111_111;
      patterns[436] = 19'b1001000100100111_111;
      patterns[437] = 19'b1010000100100111_111;
      patterns[438] = 19'b1011000100100111_111;
      patterns[439] = 19'b0100000100100000_001;
      patterns[440] = 19'b1000000100110000_000;
      patterns[441] = 19'b1001000100110000_000;
      patterns[442] = 19'b1010000100110000_000;
      patterns[443] = 19'b1011000100110000_000;
      patterns[444] = 19'b0100000100110000_001;
      patterns[445] = 19'b1000000100110001_001;
      patterns[446] = 19'b1001000100110001_001;
      patterns[447] = 19'b1010000100110001_001;
      patterns[448] = 19'b1011000100110001_001;
      patterns[449] = 19'b0100000100110000_001;
      patterns[450] = 19'b1000000100110010_010;
      patterns[451] = 19'b1001000100110010_010;
      patterns[452] = 19'b1010000100110010_010;
      patterns[453] = 19'b1011000100110010_010;
      patterns[454] = 19'b0100000100110000_001;
      patterns[455] = 19'b1000000100110011_011;
      patterns[456] = 19'b1001000100110011_011;
      patterns[457] = 19'b1010000100110011_011;
      patterns[458] = 19'b1011000100110011_011;
      patterns[459] = 19'b0100000100110000_001;
      patterns[460] = 19'b1000000100110100_100;
      patterns[461] = 19'b1001000100110100_100;
      patterns[462] = 19'b1010000100110100_100;
      patterns[463] = 19'b1011000100110100_100;
      patterns[464] = 19'b0100000100110000_001;
      patterns[465] = 19'b1000000100110101_101;
      patterns[466] = 19'b1001000100110101_101;
      patterns[467] = 19'b1010000100110101_101;
      patterns[468] = 19'b1011000100110101_101;
      patterns[469] = 19'b0100000100110000_001;
      patterns[470] = 19'b1000000100110110_110;
      patterns[471] = 19'b1001000100110110_110;
      patterns[472] = 19'b1010000100110110_110;
      patterns[473] = 19'b1011000100110110_110;
      patterns[474] = 19'b0100000100110000_001;
      patterns[475] = 19'b1000000100110111_111;
      patterns[476] = 19'b1001000100110111_111;
      patterns[477] = 19'b1010000100110111_111;
      patterns[478] = 19'b1011000100110111_111;
      patterns[479] = 19'b0100000100110000_001;
      patterns[480] = 19'b1000000101000000_000;
      patterns[481] = 19'b1001000101000000_000;
      patterns[482] = 19'b1010000101000000_000;
      patterns[483] = 19'b1011000101000000_000;
      patterns[484] = 19'b0100000101000000_001;
      patterns[485] = 19'b1000000101000001_001;
      patterns[486] = 19'b1001000101000001_001;
      patterns[487] = 19'b1010000101000001_001;
      patterns[488] = 19'b1011000101000001_001;
      patterns[489] = 19'b0100000101000000_001;
      patterns[490] = 19'b1000000101000010_010;
      patterns[491] = 19'b1001000101000010_010;
      patterns[492] = 19'b1010000101000010_010;
      patterns[493] = 19'b1011000101000010_010;
      patterns[494] = 19'b0100000101000000_001;
      patterns[495] = 19'b1000000101000011_011;
      patterns[496] = 19'b1001000101000011_011;
      patterns[497] = 19'b1010000101000011_011;
      patterns[498] = 19'b1011000101000011_011;
      patterns[499] = 19'b0100000101000000_001;
      patterns[500] = 19'b1000000101000100_100;
      patterns[501] = 19'b1001000101000100_100;
      patterns[502] = 19'b1010000101000100_100;
      patterns[503] = 19'b1011000101000100_100;
      patterns[504] = 19'b0100000101000000_001;
      patterns[505] = 19'b1000000101000101_101;
      patterns[506] = 19'b1001000101000101_101;
      patterns[507] = 19'b1010000101000101_101;
      patterns[508] = 19'b1011000101000101_101;
      patterns[509] = 19'b0100000101000000_001;
      patterns[510] = 19'b1000000101000110_110;
      patterns[511] = 19'b1001000101000110_110;
      patterns[512] = 19'b1010000101000110_110;
      patterns[513] = 19'b1011000101000110_110;
      patterns[514] = 19'b0100000101000000_001;
      patterns[515] = 19'b1000000101000111_111;
      patterns[516] = 19'b1001000101000111_111;
      patterns[517] = 19'b1010000101000111_111;
      patterns[518] = 19'b1011000101000111_111;
      patterns[519] = 19'b0100000101000000_001;
      patterns[520] = 19'b1000000101010000_000;
      patterns[521] = 19'b1001000101010000_000;
      patterns[522] = 19'b1010000101010000_000;
      patterns[523] = 19'b1011000101010000_000;
      patterns[524] = 19'b0100000101010000_001;
      patterns[525] = 19'b1000000101010001_001;
      patterns[526] = 19'b1001000101010001_001;
      patterns[527] = 19'b1010000101010001_001;
      patterns[528] = 19'b1011000101010001_001;
      patterns[529] = 19'b0100000101010000_001;
      patterns[530] = 19'b1000000101010010_010;
      patterns[531] = 19'b1001000101010010_010;
      patterns[532] = 19'b1010000101010010_010;
      patterns[533] = 19'b1011000101010010_010;
      patterns[534] = 19'b0100000101010000_001;
      patterns[535] = 19'b1000000101010011_011;
      patterns[536] = 19'b1001000101010011_011;
      patterns[537] = 19'b1010000101010011_011;
      patterns[538] = 19'b1011000101010011_011;
      patterns[539] = 19'b0100000101010000_001;
      patterns[540] = 19'b1000000101010100_100;
      patterns[541] = 19'b1001000101010100_100;
      patterns[542] = 19'b1010000101010100_100;
      patterns[543] = 19'b1011000101010100_100;
      patterns[544] = 19'b0100000101010000_001;
      patterns[545] = 19'b1000000101010101_101;
      patterns[546] = 19'b1001000101010101_101;
      patterns[547] = 19'b1010000101010101_101;
      patterns[548] = 19'b1011000101010101_101;
      patterns[549] = 19'b0100000101010000_001;
      patterns[550] = 19'b1000000101010110_110;
      patterns[551] = 19'b1001000101010110_110;
      patterns[552] = 19'b1010000101010110_110;
      patterns[553] = 19'b1011000101010110_110;
      patterns[554] = 19'b0100000101010000_001;
      patterns[555] = 19'b1000000101010111_111;
      patterns[556] = 19'b1001000101010111_111;
      patterns[557] = 19'b1010000101010111_111;
      patterns[558] = 19'b1011000101010111_111;
      patterns[559] = 19'b0100000101010000_001;
      patterns[560] = 19'b1000000101100000_000;
      patterns[561] = 19'b1001000101100000_000;
      patterns[562] = 19'b1010000101100000_000;
      patterns[563] = 19'b1011000101100000_000;
      patterns[564] = 19'b0100000101100000_001;
      patterns[565] = 19'b1000000101100001_001;
      patterns[566] = 19'b1001000101100001_001;
      patterns[567] = 19'b1010000101100001_001;
      patterns[568] = 19'b1011000101100001_001;
      patterns[569] = 19'b0100000101100000_001;
      patterns[570] = 19'b1000000101100010_010;
      patterns[571] = 19'b1001000101100010_010;
      patterns[572] = 19'b1010000101100010_010;
      patterns[573] = 19'b1011000101100010_010;
      patterns[574] = 19'b0100000101100000_001;
      patterns[575] = 19'b1000000101100011_011;
      patterns[576] = 19'b1001000101100011_011;
      patterns[577] = 19'b1010000101100011_011;
      patterns[578] = 19'b1011000101100011_011;
      patterns[579] = 19'b0100000101100000_001;
      patterns[580] = 19'b1000000101100100_100;
      patterns[581] = 19'b1001000101100100_100;
      patterns[582] = 19'b1010000101100100_100;
      patterns[583] = 19'b1011000101100100_100;
      patterns[584] = 19'b0100000101100000_001;
      patterns[585] = 19'b1000000101100101_101;
      patterns[586] = 19'b1001000101100101_101;
      patterns[587] = 19'b1010000101100101_101;
      patterns[588] = 19'b1011000101100101_101;
      patterns[589] = 19'b0100000101100000_001;
      patterns[590] = 19'b1000000101100110_110;
      patterns[591] = 19'b1001000101100110_110;
      patterns[592] = 19'b1010000101100110_110;
      patterns[593] = 19'b1011000101100110_110;
      patterns[594] = 19'b0100000101100000_001;
      patterns[595] = 19'b1000000101100111_111;
      patterns[596] = 19'b1001000101100111_111;
      patterns[597] = 19'b1010000101100111_111;
      patterns[598] = 19'b1011000101100111_111;
      patterns[599] = 19'b0100000101100000_001;
      patterns[600] = 19'b1000000101110000_000;
      patterns[601] = 19'b1001000101110000_000;
      patterns[602] = 19'b1010000101110000_000;
      patterns[603] = 19'b1011000101110000_000;
      patterns[604] = 19'b0100000101110000_001;
      patterns[605] = 19'b1000000101110001_001;
      patterns[606] = 19'b1001000101110001_001;
      patterns[607] = 19'b1010000101110001_001;
      patterns[608] = 19'b1011000101110001_001;
      patterns[609] = 19'b0100000101110000_001;
      patterns[610] = 19'b1000000101110010_010;
      patterns[611] = 19'b1001000101110010_010;
      patterns[612] = 19'b1010000101110010_010;
      patterns[613] = 19'b1011000101110010_010;
      patterns[614] = 19'b0100000101110000_001;
      patterns[615] = 19'b1000000101110011_011;
      patterns[616] = 19'b1001000101110011_011;
      patterns[617] = 19'b1010000101110011_011;
      patterns[618] = 19'b1011000101110011_011;
      patterns[619] = 19'b0100000101110000_001;
      patterns[620] = 19'b1000000101110100_100;
      patterns[621] = 19'b1001000101110100_100;
      patterns[622] = 19'b1010000101110100_100;
      patterns[623] = 19'b1011000101110100_100;
      patterns[624] = 19'b0100000101110000_001;
      patterns[625] = 19'b1000000101110101_101;
      patterns[626] = 19'b1001000101110101_101;
      patterns[627] = 19'b1010000101110101_101;
      patterns[628] = 19'b1011000101110101_101;
      patterns[629] = 19'b0100000101110000_001;
      patterns[630] = 19'b1000000101110110_110;
      patterns[631] = 19'b1001000101110110_110;
      patterns[632] = 19'b1010000101110110_110;
      patterns[633] = 19'b1011000101110110_110;
      patterns[634] = 19'b0100000101110000_001;
      patterns[635] = 19'b1000000101110111_111;
      patterns[636] = 19'b1001000101110111_111;
      patterns[637] = 19'b1010000101110111_111;
      patterns[638] = 19'b1011000101110111_111;
      patterns[639] = 19'b0100000101110000_001;
      patterns[640] = 19'b1000001000000000_000;
      patterns[641] = 19'b1001001000000000_000;
      patterns[642] = 19'b1010001000000000_000;
      patterns[643] = 19'b1011001000000000_000;
      patterns[644] = 19'b0100001000000000_010;
      patterns[645] = 19'b1000001000000001_001;
      patterns[646] = 19'b1001001000000001_001;
      patterns[647] = 19'b1010001000000001_001;
      patterns[648] = 19'b1011001000000001_001;
      patterns[649] = 19'b0100001000000000_010;
      patterns[650] = 19'b1000001000000010_010;
      patterns[651] = 19'b1001001000000010_010;
      patterns[652] = 19'b1010001000000010_010;
      patterns[653] = 19'b1011001000000010_010;
      patterns[654] = 19'b0100001000000000_010;
      patterns[655] = 19'b1000001000000011_011;
      patterns[656] = 19'b1001001000000011_011;
      patterns[657] = 19'b1010001000000011_011;
      patterns[658] = 19'b1011001000000011_011;
      patterns[659] = 19'b0100001000000000_010;
      patterns[660] = 19'b1000001000000100_100;
      patterns[661] = 19'b1001001000000100_100;
      patterns[662] = 19'b1010001000000100_100;
      patterns[663] = 19'b1011001000000100_100;
      patterns[664] = 19'b0100001000000000_010;
      patterns[665] = 19'b1000001000000101_101;
      patterns[666] = 19'b1001001000000101_101;
      patterns[667] = 19'b1010001000000101_101;
      patterns[668] = 19'b1011001000000101_101;
      patterns[669] = 19'b0100001000000000_010;
      patterns[670] = 19'b1000001000000110_110;
      patterns[671] = 19'b1001001000000110_110;
      patterns[672] = 19'b1010001000000110_110;
      patterns[673] = 19'b1011001000000110_110;
      patterns[674] = 19'b0100001000000000_010;
      patterns[675] = 19'b1000001000000111_111;
      patterns[676] = 19'b1001001000000111_111;
      patterns[677] = 19'b1010001000000111_111;
      patterns[678] = 19'b1011001000000111_111;
      patterns[679] = 19'b0100001000000000_010;
      patterns[680] = 19'b1000001000010000_000;
      patterns[681] = 19'b1001001000010000_000;
      patterns[682] = 19'b1010001000010000_000;
      patterns[683] = 19'b1011001000010000_000;
      patterns[684] = 19'b0100001000010000_010;
      patterns[685] = 19'b1000001000010001_001;
      patterns[686] = 19'b1001001000010001_001;
      patterns[687] = 19'b1010001000010001_001;
      patterns[688] = 19'b1011001000010001_001;
      patterns[689] = 19'b0100001000010000_010;
      patterns[690] = 19'b1000001000010010_010;
      patterns[691] = 19'b1001001000010010_010;
      patterns[692] = 19'b1010001000010010_010;
      patterns[693] = 19'b1011001000010010_010;
      patterns[694] = 19'b0100001000010000_010;
      patterns[695] = 19'b1000001000010011_011;
      patterns[696] = 19'b1001001000010011_011;
      patterns[697] = 19'b1010001000010011_011;
      patterns[698] = 19'b1011001000010011_011;
      patterns[699] = 19'b0100001000010000_010;
      patterns[700] = 19'b1000001000010100_100;
      patterns[701] = 19'b1001001000010100_100;
      patterns[702] = 19'b1010001000010100_100;
      patterns[703] = 19'b1011001000010100_100;
      patterns[704] = 19'b0100001000010000_010;
      patterns[705] = 19'b1000001000010101_101;
      patterns[706] = 19'b1001001000010101_101;
      patterns[707] = 19'b1010001000010101_101;
      patterns[708] = 19'b1011001000010101_101;
      patterns[709] = 19'b0100001000010000_010;
      patterns[710] = 19'b1000001000010110_110;
      patterns[711] = 19'b1001001000010110_110;
      patterns[712] = 19'b1010001000010110_110;
      patterns[713] = 19'b1011001000010110_110;
      patterns[714] = 19'b0100001000010000_010;
      patterns[715] = 19'b1000001000010111_111;
      patterns[716] = 19'b1001001000010111_111;
      patterns[717] = 19'b1010001000010111_111;
      patterns[718] = 19'b1011001000010111_111;
      patterns[719] = 19'b0100001000010000_010;
      patterns[720] = 19'b1000001000100000_000;
      patterns[721] = 19'b1001001000100000_000;
      patterns[722] = 19'b1010001000100000_000;
      patterns[723] = 19'b1011001000100000_000;
      patterns[724] = 19'b0100001000100000_010;
      patterns[725] = 19'b1000001000100001_001;
      patterns[726] = 19'b1001001000100001_001;
      patterns[727] = 19'b1010001000100001_001;
      patterns[728] = 19'b1011001000100001_001;
      patterns[729] = 19'b0100001000100000_010;
      patterns[730] = 19'b1000001000100010_010;
      patterns[731] = 19'b1001001000100010_010;
      patterns[732] = 19'b1010001000100010_010;
      patterns[733] = 19'b1011001000100010_010;
      patterns[734] = 19'b0100001000100000_010;
      patterns[735] = 19'b1000001000100011_011;
      patterns[736] = 19'b1001001000100011_011;
      patterns[737] = 19'b1010001000100011_011;
      patterns[738] = 19'b1011001000100011_011;
      patterns[739] = 19'b0100001000100000_010;
      patterns[740] = 19'b1000001000100100_100;
      patterns[741] = 19'b1001001000100100_100;
      patterns[742] = 19'b1010001000100100_100;
      patterns[743] = 19'b1011001000100100_100;
      patterns[744] = 19'b0100001000100000_010;
      patterns[745] = 19'b1000001000100101_101;
      patterns[746] = 19'b1001001000100101_101;
      patterns[747] = 19'b1010001000100101_101;
      patterns[748] = 19'b1011001000100101_101;
      patterns[749] = 19'b0100001000100000_010;
      patterns[750] = 19'b1000001000100110_110;
      patterns[751] = 19'b1001001000100110_110;
      patterns[752] = 19'b1010001000100110_110;
      patterns[753] = 19'b1011001000100110_110;
      patterns[754] = 19'b0100001000100000_010;
      patterns[755] = 19'b1000001000100111_111;
      patterns[756] = 19'b1001001000100111_111;
      patterns[757] = 19'b1010001000100111_111;
      patterns[758] = 19'b1011001000100111_111;
      patterns[759] = 19'b0100001000100000_010;
      patterns[760] = 19'b1000001000110000_000;
      patterns[761] = 19'b1001001000110000_000;
      patterns[762] = 19'b1010001000110000_000;
      patterns[763] = 19'b1011001000110000_000;
      patterns[764] = 19'b0100001000110000_010;
      patterns[765] = 19'b1000001000110001_001;
      patterns[766] = 19'b1001001000110001_001;
      patterns[767] = 19'b1010001000110001_001;
      patterns[768] = 19'b1011001000110001_001;
      patterns[769] = 19'b0100001000110000_010;
      patterns[770] = 19'b1000001000110010_010;
      patterns[771] = 19'b1001001000110010_010;
      patterns[772] = 19'b1010001000110010_010;
      patterns[773] = 19'b1011001000110010_010;
      patterns[774] = 19'b0100001000110000_010;
      patterns[775] = 19'b1000001000110011_011;
      patterns[776] = 19'b1001001000110011_011;
      patterns[777] = 19'b1010001000110011_011;
      patterns[778] = 19'b1011001000110011_011;
      patterns[779] = 19'b0100001000110000_010;
      patterns[780] = 19'b1000001000110100_100;
      patterns[781] = 19'b1001001000110100_100;
      patterns[782] = 19'b1010001000110100_100;
      patterns[783] = 19'b1011001000110100_100;
      patterns[784] = 19'b0100001000110000_010;
      patterns[785] = 19'b1000001000110101_101;
      patterns[786] = 19'b1001001000110101_101;
      patterns[787] = 19'b1010001000110101_101;
      patterns[788] = 19'b1011001000110101_101;
      patterns[789] = 19'b0100001000110000_010;
      patterns[790] = 19'b1000001000110110_110;
      patterns[791] = 19'b1001001000110110_110;
      patterns[792] = 19'b1010001000110110_110;
      patterns[793] = 19'b1011001000110110_110;
      patterns[794] = 19'b0100001000110000_010;
      patterns[795] = 19'b1000001000110111_111;
      patterns[796] = 19'b1001001000110111_111;
      patterns[797] = 19'b1010001000110111_111;
      patterns[798] = 19'b1011001000110111_111;
      patterns[799] = 19'b0100001000110000_010;
      patterns[800] = 19'b1000001001000000_000;
      patterns[801] = 19'b1001001001000000_000;
      patterns[802] = 19'b1010001001000000_000;
      patterns[803] = 19'b1011001001000000_000;
      patterns[804] = 19'b0100001001000000_010;
      patterns[805] = 19'b1000001001000001_001;
      patterns[806] = 19'b1001001001000001_001;
      patterns[807] = 19'b1010001001000001_001;
      patterns[808] = 19'b1011001001000001_001;
      patterns[809] = 19'b0100001001000000_010;
      patterns[810] = 19'b1000001001000010_010;
      patterns[811] = 19'b1001001001000010_010;
      patterns[812] = 19'b1010001001000010_010;
      patterns[813] = 19'b1011001001000010_010;
      patterns[814] = 19'b0100001001000000_010;
      patterns[815] = 19'b1000001001000011_011;
      patterns[816] = 19'b1001001001000011_011;
      patterns[817] = 19'b1010001001000011_011;
      patterns[818] = 19'b1011001001000011_011;
      patterns[819] = 19'b0100001001000000_010;
      patterns[820] = 19'b1000001001000100_100;
      patterns[821] = 19'b1001001001000100_100;
      patterns[822] = 19'b1010001001000100_100;
      patterns[823] = 19'b1011001001000100_100;
      patterns[824] = 19'b0100001001000000_010;
      patterns[825] = 19'b1000001001000101_101;
      patterns[826] = 19'b1001001001000101_101;
      patterns[827] = 19'b1010001001000101_101;
      patterns[828] = 19'b1011001001000101_101;
      patterns[829] = 19'b0100001001000000_010;
      patterns[830] = 19'b1000001001000110_110;
      patterns[831] = 19'b1001001001000110_110;
      patterns[832] = 19'b1010001001000110_110;
      patterns[833] = 19'b1011001001000110_110;
      patterns[834] = 19'b0100001001000000_010;
      patterns[835] = 19'b1000001001000111_111;
      patterns[836] = 19'b1001001001000111_111;
      patterns[837] = 19'b1010001001000111_111;
      patterns[838] = 19'b1011001001000111_111;
      patterns[839] = 19'b0100001001000000_010;
      patterns[840] = 19'b1000001001010000_000;
      patterns[841] = 19'b1001001001010000_000;
      patterns[842] = 19'b1010001001010000_000;
      patterns[843] = 19'b1011001001010000_000;
      patterns[844] = 19'b0100001001010000_010;
      patterns[845] = 19'b1000001001010001_001;
      patterns[846] = 19'b1001001001010001_001;
      patterns[847] = 19'b1010001001010001_001;
      patterns[848] = 19'b1011001001010001_001;
      patterns[849] = 19'b0100001001010000_010;
      patterns[850] = 19'b1000001001010010_010;
      patterns[851] = 19'b1001001001010010_010;
      patterns[852] = 19'b1010001001010010_010;
      patterns[853] = 19'b1011001001010010_010;
      patterns[854] = 19'b0100001001010000_010;
      patterns[855] = 19'b1000001001010011_011;
      patterns[856] = 19'b1001001001010011_011;
      patterns[857] = 19'b1010001001010011_011;
      patterns[858] = 19'b1011001001010011_011;
      patterns[859] = 19'b0100001001010000_010;
      patterns[860] = 19'b1000001001010100_100;
      patterns[861] = 19'b1001001001010100_100;
      patterns[862] = 19'b1010001001010100_100;
      patterns[863] = 19'b1011001001010100_100;
      patterns[864] = 19'b0100001001010000_010;
      patterns[865] = 19'b1000001001010101_101;
      patterns[866] = 19'b1001001001010101_101;
      patterns[867] = 19'b1010001001010101_101;
      patterns[868] = 19'b1011001001010101_101;
      patterns[869] = 19'b0100001001010000_010;
      patterns[870] = 19'b1000001001010110_110;
      patterns[871] = 19'b1001001001010110_110;
      patterns[872] = 19'b1010001001010110_110;
      patterns[873] = 19'b1011001001010110_110;
      patterns[874] = 19'b0100001001010000_010;
      patterns[875] = 19'b1000001001010111_111;
      patterns[876] = 19'b1001001001010111_111;
      patterns[877] = 19'b1010001001010111_111;
      patterns[878] = 19'b1011001001010111_111;
      patterns[879] = 19'b0100001001010000_010;
      patterns[880] = 19'b1000001001100000_000;
      patterns[881] = 19'b1001001001100000_000;
      patterns[882] = 19'b1010001001100000_000;
      patterns[883] = 19'b1011001001100000_000;
      patterns[884] = 19'b0100001001100000_010;
      patterns[885] = 19'b1000001001100001_001;
      patterns[886] = 19'b1001001001100001_001;
      patterns[887] = 19'b1010001001100001_001;
      patterns[888] = 19'b1011001001100001_001;
      patterns[889] = 19'b0100001001100000_010;
      patterns[890] = 19'b1000001001100010_010;
      patterns[891] = 19'b1001001001100010_010;
      patterns[892] = 19'b1010001001100010_010;
      patterns[893] = 19'b1011001001100010_010;
      patterns[894] = 19'b0100001001100000_010;
      patterns[895] = 19'b1000001001100011_011;
      patterns[896] = 19'b1001001001100011_011;
      patterns[897] = 19'b1010001001100011_011;
      patterns[898] = 19'b1011001001100011_011;
      patterns[899] = 19'b0100001001100000_010;
      patterns[900] = 19'b1000001001100100_100;
      patterns[901] = 19'b1001001001100100_100;
      patterns[902] = 19'b1010001001100100_100;
      patterns[903] = 19'b1011001001100100_100;
      patterns[904] = 19'b0100001001100000_010;
      patterns[905] = 19'b1000001001100101_101;
      patterns[906] = 19'b1001001001100101_101;
      patterns[907] = 19'b1010001001100101_101;
      patterns[908] = 19'b1011001001100101_101;
      patterns[909] = 19'b0100001001100000_010;
      patterns[910] = 19'b1000001001100110_110;
      patterns[911] = 19'b1001001001100110_110;
      patterns[912] = 19'b1010001001100110_110;
      patterns[913] = 19'b1011001001100110_110;
      patterns[914] = 19'b0100001001100000_010;
      patterns[915] = 19'b1000001001100111_111;
      patterns[916] = 19'b1001001001100111_111;
      patterns[917] = 19'b1010001001100111_111;
      patterns[918] = 19'b1011001001100111_111;
      patterns[919] = 19'b0100001001100000_010;
      patterns[920] = 19'b1000001001110000_000;
      patterns[921] = 19'b1001001001110000_000;
      patterns[922] = 19'b1010001001110000_000;
      patterns[923] = 19'b1011001001110000_000;
      patterns[924] = 19'b0100001001110000_010;
      patterns[925] = 19'b1000001001110001_001;
      patterns[926] = 19'b1001001001110001_001;
      patterns[927] = 19'b1010001001110001_001;
      patterns[928] = 19'b1011001001110001_001;
      patterns[929] = 19'b0100001001110000_010;
      patterns[930] = 19'b1000001001110010_010;
      patterns[931] = 19'b1001001001110010_010;
      patterns[932] = 19'b1010001001110010_010;
      patterns[933] = 19'b1011001001110010_010;
      patterns[934] = 19'b0100001001110000_010;
      patterns[935] = 19'b1000001001110011_011;
      patterns[936] = 19'b1001001001110011_011;
      patterns[937] = 19'b1010001001110011_011;
      patterns[938] = 19'b1011001001110011_011;
      patterns[939] = 19'b0100001001110000_010;
      patterns[940] = 19'b1000001001110100_100;
      patterns[941] = 19'b1001001001110100_100;
      patterns[942] = 19'b1010001001110100_100;
      patterns[943] = 19'b1011001001110100_100;
      patterns[944] = 19'b0100001001110000_010;
      patterns[945] = 19'b1000001001110101_101;
      patterns[946] = 19'b1001001001110101_101;
      patterns[947] = 19'b1010001001110101_101;
      patterns[948] = 19'b1011001001110101_101;
      patterns[949] = 19'b0100001001110000_010;
      patterns[950] = 19'b1000001001110110_110;
      patterns[951] = 19'b1001001001110110_110;
      patterns[952] = 19'b1010001001110110_110;
      patterns[953] = 19'b1011001001110110_110;
      patterns[954] = 19'b0100001001110000_010;
      patterns[955] = 19'b1000001001110111_111;
      patterns[956] = 19'b1001001001110111_111;
      patterns[957] = 19'b1010001001110111_111;
      patterns[958] = 19'b1011001001110111_111;
      patterns[959] = 19'b0100001001110000_010;
      patterns[960] = 19'b1000001100000000_000;
      patterns[961] = 19'b1001001100000000_000;
      patterns[962] = 19'b1010001100000000_000;
      patterns[963] = 19'b1011001100000000_000;
      patterns[964] = 19'b0100001100000000_011;
      patterns[965] = 19'b1000001100000001_001;
      patterns[966] = 19'b1001001100000001_001;
      patterns[967] = 19'b1010001100000001_001;
      patterns[968] = 19'b1011001100000001_001;
      patterns[969] = 19'b0100001100000000_011;
      patterns[970] = 19'b1000001100000010_010;
      patterns[971] = 19'b1001001100000010_010;
      patterns[972] = 19'b1010001100000010_010;
      patterns[973] = 19'b1011001100000010_010;
      patterns[974] = 19'b0100001100000000_011;
      patterns[975] = 19'b1000001100000011_011;
      patterns[976] = 19'b1001001100000011_011;
      patterns[977] = 19'b1010001100000011_011;
      patterns[978] = 19'b1011001100000011_011;
      patterns[979] = 19'b0100001100000000_011;
      patterns[980] = 19'b1000001100000100_100;
      patterns[981] = 19'b1001001100000100_100;
      patterns[982] = 19'b1010001100000100_100;
      patterns[983] = 19'b1011001100000100_100;
      patterns[984] = 19'b0100001100000000_011;
      patterns[985] = 19'b1000001100000101_101;
      patterns[986] = 19'b1001001100000101_101;
      patterns[987] = 19'b1010001100000101_101;
      patterns[988] = 19'b1011001100000101_101;
      patterns[989] = 19'b0100001100000000_011;
      patterns[990] = 19'b1000001100000110_110;
      patterns[991] = 19'b1001001100000110_110;
      patterns[992] = 19'b1010001100000110_110;
      patterns[993] = 19'b1011001100000110_110;
      patterns[994] = 19'b0100001100000000_011;
      patterns[995] = 19'b1000001100000111_111;
      patterns[996] = 19'b1001001100000111_111;
      patterns[997] = 19'b1010001100000111_111;
      patterns[998] = 19'b1011001100000111_111;
      patterns[999] = 19'b0100001100000000_011;
      patterns[1000] = 19'b1000001100010000_000;
      patterns[1001] = 19'b1001001100010000_000;
      patterns[1002] = 19'b1010001100010000_000;
      patterns[1003] = 19'b1011001100010000_000;
      patterns[1004] = 19'b0100001100010000_011;
      patterns[1005] = 19'b1000001100010001_001;
      patterns[1006] = 19'b1001001100010001_001;
      patterns[1007] = 19'b1010001100010001_001;
      patterns[1008] = 19'b1011001100010001_001;
      patterns[1009] = 19'b0100001100010000_011;
      patterns[1010] = 19'b1000001100010010_010;
      patterns[1011] = 19'b1001001100010010_010;
      patterns[1012] = 19'b1010001100010010_010;
      patterns[1013] = 19'b1011001100010010_010;
      patterns[1014] = 19'b0100001100010000_011;
      patterns[1015] = 19'b1000001100010011_011;
      patterns[1016] = 19'b1001001100010011_011;
      patterns[1017] = 19'b1010001100010011_011;
      patterns[1018] = 19'b1011001100010011_011;
      patterns[1019] = 19'b0100001100010000_011;
      patterns[1020] = 19'b1000001100010100_100;
      patterns[1021] = 19'b1001001100010100_100;
      patterns[1022] = 19'b1010001100010100_100;
      patterns[1023] = 19'b1011001100010100_100;
      patterns[1024] = 19'b0100001100010000_011;
      patterns[1025] = 19'b1000001100010101_101;
      patterns[1026] = 19'b1001001100010101_101;
      patterns[1027] = 19'b1010001100010101_101;
      patterns[1028] = 19'b1011001100010101_101;
      patterns[1029] = 19'b0100001100010000_011;
      patterns[1030] = 19'b1000001100010110_110;
      patterns[1031] = 19'b1001001100010110_110;
      patterns[1032] = 19'b1010001100010110_110;
      patterns[1033] = 19'b1011001100010110_110;
      patterns[1034] = 19'b0100001100010000_011;
      patterns[1035] = 19'b1000001100010111_111;
      patterns[1036] = 19'b1001001100010111_111;
      patterns[1037] = 19'b1010001100010111_111;
      patterns[1038] = 19'b1011001100010111_111;
      patterns[1039] = 19'b0100001100010000_011;
      patterns[1040] = 19'b1000001100100000_000;
      patterns[1041] = 19'b1001001100100000_000;
      patterns[1042] = 19'b1010001100100000_000;
      patterns[1043] = 19'b1011001100100000_000;
      patterns[1044] = 19'b0100001100100000_011;
      patterns[1045] = 19'b1000001100100001_001;
      patterns[1046] = 19'b1001001100100001_001;
      patterns[1047] = 19'b1010001100100001_001;
      patterns[1048] = 19'b1011001100100001_001;
      patterns[1049] = 19'b0100001100100000_011;
      patterns[1050] = 19'b1000001100100010_010;
      patterns[1051] = 19'b1001001100100010_010;
      patterns[1052] = 19'b1010001100100010_010;
      patterns[1053] = 19'b1011001100100010_010;
      patterns[1054] = 19'b0100001100100000_011;
      patterns[1055] = 19'b1000001100100011_011;
      patterns[1056] = 19'b1001001100100011_011;
      patterns[1057] = 19'b1010001100100011_011;
      patterns[1058] = 19'b1011001100100011_011;
      patterns[1059] = 19'b0100001100100000_011;
      patterns[1060] = 19'b1000001100100100_100;
      patterns[1061] = 19'b1001001100100100_100;
      patterns[1062] = 19'b1010001100100100_100;
      patterns[1063] = 19'b1011001100100100_100;
      patterns[1064] = 19'b0100001100100000_011;
      patterns[1065] = 19'b1000001100100101_101;
      patterns[1066] = 19'b1001001100100101_101;
      patterns[1067] = 19'b1010001100100101_101;
      patterns[1068] = 19'b1011001100100101_101;
      patterns[1069] = 19'b0100001100100000_011;
      patterns[1070] = 19'b1000001100100110_110;
      patterns[1071] = 19'b1001001100100110_110;
      patterns[1072] = 19'b1010001100100110_110;
      patterns[1073] = 19'b1011001100100110_110;
      patterns[1074] = 19'b0100001100100000_011;
      patterns[1075] = 19'b1000001100100111_111;
      patterns[1076] = 19'b1001001100100111_111;
      patterns[1077] = 19'b1010001100100111_111;
      patterns[1078] = 19'b1011001100100111_111;
      patterns[1079] = 19'b0100001100100000_011;
      patterns[1080] = 19'b1000001100110000_000;
      patterns[1081] = 19'b1001001100110000_000;
      patterns[1082] = 19'b1010001100110000_000;
      patterns[1083] = 19'b1011001100110000_000;
      patterns[1084] = 19'b0100001100110000_011;
      patterns[1085] = 19'b1000001100110001_001;
      patterns[1086] = 19'b1001001100110001_001;
      patterns[1087] = 19'b1010001100110001_001;
      patterns[1088] = 19'b1011001100110001_001;
      patterns[1089] = 19'b0100001100110000_011;
      patterns[1090] = 19'b1000001100110010_010;
      patterns[1091] = 19'b1001001100110010_010;
      patterns[1092] = 19'b1010001100110010_010;
      patterns[1093] = 19'b1011001100110010_010;
      patterns[1094] = 19'b0100001100110000_011;
      patterns[1095] = 19'b1000001100110011_011;
      patterns[1096] = 19'b1001001100110011_011;
      patterns[1097] = 19'b1010001100110011_011;
      patterns[1098] = 19'b1011001100110011_011;
      patterns[1099] = 19'b0100001100110000_011;
      patterns[1100] = 19'b1000001100110100_100;
      patterns[1101] = 19'b1001001100110100_100;
      patterns[1102] = 19'b1010001100110100_100;
      patterns[1103] = 19'b1011001100110100_100;
      patterns[1104] = 19'b0100001100110000_011;
      patterns[1105] = 19'b1000001100110101_101;
      patterns[1106] = 19'b1001001100110101_101;
      patterns[1107] = 19'b1010001100110101_101;
      patterns[1108] = 19'b1011001100110101_101;
      patterns[1109] = 19'b0100001100110000_011;
      patterns[1110] = 19'b1000001100110110_110;
      patterns[1111] = 19'b1001001100110110_110;
      patterns[1112] = 19'b1010001100110110_110;
      patterns[1113] = 19'b1011001100110110_110;
      patterns[1114] = 19'b0100001100110000_011;
      patterns[1115] = 19'b1000001100110111_111;
      patterns[1116] = 19'b1001001100110111_111;
      patterns[1117] = 19'b1010001100110111_111;
      patterns[1118] = 19'b1011001100110111_111;
      patterns[1119] = 19'b0100001100110000_011;
      patterns[1120] = 19'b1000001101000000_000;
      patterns[1121] = 19'b1001001101000000_000;
      patterns[1122] = 19'b1010001101000000_000;
      patterns[1123] = 19'b1011001101000000_000;
      patterns[1124] = 19'b0100001101000000_011;
      patterns[1125] = 19'b1000001101000001_001;
      patterns[1126] = 19'b1001001101000001_001;
      patterns[1127] = 19'b1010001101000001_001;
      patterns[1128] = 19'b1011001101000001_001;
      patterns[1129] = 19'b0100001101000000_011;
      patterns[1130] = 19'b1000001101000010_010;
      patterns[1131] = 19'b1001001101000010_010;
      patterns[1132] = 19'b1010001101000010_010;
      patterns[1133] = 19'b1011001101000010_010;
      patterns[1134] = 19'b0100001101000000_011;
      patterns[1135] = 19'b1000001101000011_011;
      patterns[1136] = 19'b1001001101000011_011;
      patterns[1137] = 19'b1010001101000011_011;
      patterns[1138] = 19'b1011001101000011_011;
      patterns[1139] = 19'b0100001101000000_011;
      patterns[1140] = 19'b1000001101000100_100;
      patterns[1141] = 19'b1001001101000100_100;
      patterns[1142] = 19'b1010001101000100_100;
      patterns[1143] = 19'b1011001101000100_100;
      patterns[1144] = 19'b0100001101000000_011;
      patterns[1145] = 19'b1000001101000101_101;
      patterns[1146] = 19'b1001001101000101_101;
      patterns[1147] = 19'b1010001101000101_101;
      patterns[1148] = 19'b1011001101000101_101;
      patterns[1149] = 19'b0100001101000000_011;
      patterns[1150] = 19'b1000001101000110_110;
      patterns[1151] = 19'b1001001101000110_110;
      patterns[1152] = 19'b1010001101000110_110;
      patterns[1153] = 19'b1011001101000110_110;
      patterns[1154] = 19'b0100001101000000_011;
      patterns[1155] = 19'b1000001101000111_111;
      patterns[1156] = 19'b1001001101000111_111;
      patterns[1157] = 19'b1010001101000111_111;
      patterns[1158] = 19'b1011001101000111_111;
      patterns[1159] = 19'b0100001101000000_011;
      patterns[1160] = 19'b1000001101010000_000;
      patterns[1161] = 19'b1001001101010000_000;
      patterns[1162] = 19'b1010001101010000_000;
      patterns[1163] = 19'b1011001101010000_000;
      patterns[1164] = 19'b0100001101010000_011;
      patterns[1165] = 19'b1000001101010001_001;
      patterns[1166] = 19'b1001001101010001_001;
      patterns[1167] = 19'b1010001101010001_001;
      patterns[1168] = 19'b1011001101010001_001;
      patterns[1169] = 19'b0100001101010000_011;
      patterns[1170] = 19'b1000001101010010_010;
      patterns[1171] = 19'b1001001101010010_010;
      patterns[1172] = 19'b1010001101010010_010;
      patterns[1173] = 19'b1011001101010010_010;
      patterns[1174] = 19'b0100001101010000_011;
      patterns[1175] = 19'b1000001101010011_011;
      patterns[1176] = 19'b1001001101010011_011;
      patterns[1177] = 19'b1010001101010011_011;
      patterns[1178] = 19'b1011001101010011_011;
      patterns[1179] = 19'b0100001101010000_011;
      patterns[1180] = 19'b1000001101010100_100;
      patterns[1181] = 19'b1001001101010100_100;
      patterns[1182] = 19'b1010001101010100_100;
      patterns[1183] = 19'b1011001101010100_100;
      patterns[1184] = 19'b0100001101010000_011;
      patterns[1185] = 19'b1000001101010101_101;
      patterns[1186] = 19'b1001001101010101_101;
      patterns[1187] = 19'b1010001101010101_101;
      patterns[1188] = 19'b1011001101010101_101;
      patterns[1189] = 19'b0100001101010000_011;
      patterns[1190] = 19'b1000001101010110_110;
      patterns[1191] = 19'b1001001101010110_110;
      patterns[1192] = 19'b1010001101010110_110;
      patterns[1193] = 19'b1011001101010110_110;
      patterns[1194] = 19'b0100001101010000_011;
      patterns[1195] = 19'b1000001101010111_111;
      patterns[1196] = 19'b1001001101010111_111;
      patterns[1197] = 19'b1010001101010111_111;
      patterns[1198] = 19'b1011001101010111_111;
      patterns[1199] = 19'b0100001101010000_011;
      patterns[1200] = 19'b1000001101100000_000;
      patterns[1201] = 19'b1001001101100000_000;
      patterns[1202] = 19'b1010001101100000_000;
      patterns[1203] = 19'b1011001101100000_000;
      patterns[1204] = 19'b0100001101100000_011;
      patterns[1205] = 19'b1000001101100001_001;
      patterns[1206] = 19'b1001001101100001_001;
      patterns[1207] = 19'b1010001101100001_001;
      patterns[1208] = 19'b1011001101100001_001;
      patterns[1209] = 19'b0100001101100000_011;
      patterns[1210] = 19'b1000001101100010_010;
      patterns[1211] = 19'b1001001101100010_010;
      patterns[1212] = 19'b1010001101100010_010;
      patterns[1213] = 19'b1011001101100010_010;
      patterns[1214] = 19'b0100001101100000_011;
      patterns[1215] = 19'b1000001101100011_011;
      patterns[1216] = 19'b1001001101100011_011;
      patterns[1217] = 19'b1010001101100011_011;
      patterns[1218] = 19'b1011001101100011_011;
      patterns[1219] = 19'b0100001101100000_011;
      patterns[1220] = 19'b1000001101100100_100;
      patterns[1221] = 19'b1001001101100100_100;
      patterns[1222] = 19'b1010001101100100_100;
      patterns[1223] = 19'b1011001101100100_100;
      patterns[1224] = 19'b0100001101100000_011;
      patterns[1225] = 19'b1000001101100101_101;
      patterns[1226] = 19'b1001001101100101_101;
      patterns[1227] = 19'b1010001101100101_101;
      patterns[1228] = 19'b1011001101100101_101;
      patterns[1229] = 19'b0100001101100000_011;
      patterns[1230] = 19'b1000001101100110_110;
      patterns[1231] = 19'b1001001101100110_110;
      patterns[1232] = 19'b1010001101100110_110;
      patterns[1233] = 19'b1011001101100110_110;
      patterns[1234] = 19'b0100001101100000_011;
      patterns[1235] = 19'b1000001101100111_111;
      patterns[1236] = 19'b1001001101100111_111;
      patterns[1237] = 19'b1010001101100111_111;
      patterns[1238] = 19'b1011001101100111_111;
      patterns[1239] = 19'b0100001101100000_011;
      patterns[1240] = 19'b1000001101110000_000;
      patterns[1241] = 19'b1001001101110000_000;
      patterns[1242] = 19'b1010001101110000_000;
      patterns[1243] = 19'b1011001101110000_000;
      patterns[1244] = 19'b0100001101110000_011;
      patterns[1245] = 19'b1000001101110001_001;
      patterns[1246] = 19'b1001001101110001_001;
      patterns[1247] = 19'b1010001101110001_001;
      patterns[1248] = 19'b1011001101110001_001;
      patterns[1249] = 19'b0100001101110000_011;
      patterns[1250] = 19'b1000001101110010_010;
      patterns[1251] = 19'b1001001101110010_010;
      patterns[1252] = 19'b1010001101110010_010;
      patterns[1253] = 19'b1011001101110010_010;
      patterns[1254] = 19'b0100001101110000_011;
      patterns[1255] = 19'b1000001101110011_011;
      patterns[1256] = 19'b1001001101110011_011;
      patterns[1257] = 19'b1010001101110011_011;
      patterns[1258] = 19'b1011001101110011_011;
      patterns[1259] = 19'b0100001101110000_011;
      patterns[1260] = 19'b1000001101110100_100;
      patterns[1261] = 19'b1001001101110100_100;
      patterns[1262] = 19'b1010001101110100_100;
      patterns[1263] = 19'b1011001101110100_100;
      patterns[1264] = 19'b0100001101110000_011;
      patterns[1265] = 19'b1000001101110101_101;
      patterns[1266] = 19'b1001001101110101_101;
      patterns[1267] = 19'b1010001101110101_101;
      patterns[1268] = 19'b1011001101110101_101;
      patterns[1269] = 19'b0100001101110000_011;
      patterns[1270] = 19'b1000001101110110_110;
      patterns[1271] = 19'b1001001101110110_110;
      patterns[1272] = 19'b1010001101110110_110;
      patterns[1273] = 19'b1011001101110110_110;
      patterns[1274] = 19'b0100001101110000_011;
      patterns[1275] = 19'b1000001101110111_111;
      patterns[1276] = 19'b1001001101110111_111;
      patterns[1277] = 19'b1010001101110111_111;
      patterns[1278] = 19'b1011001101110111_111;
      patterns[1279] = 19'b0100001101110000_011;
      patterns[1280] = 19'b1000010000000000_000;
      patterns[1281] = 19'b1001010000000000_000;
      patterns[1282] = 19'b1010010000000000_000;
      patterns[1283] = 19'b1011010000000000_000;
      patterns[1284] = 19'b0100010000000000_100;
      patterns[1285] = 19'b1000010000000001_001;
      patterns[1286] = 19'b1001010000000001_001;
      patterns[1287] = 19'b1010010000000001_001;
      patterns[1288] = 19'b1011010000000001_001;
      patterns[1289] = 19'b0100010000000000_100;
      patterns[1290] = 19'b1000010000000010_010;
      patterns[1291] = 19'b1001010000000010_010;
      patterns[1292] = 19'b1010010000000010_010;
      patterns[1293] = 19'b1011010000000010_010;
      patterns[1294] = 19'b0100010000000000_100;
      patterns[1295] = 19'b1000010000000011_011;
      patterns[1296] = 19'b1001010000000011_011;
      patterns[1297] = 19'b1010010000000011_011;
      patterns[1298] = 19'b1011010000000011_011;
      patterns[1299] = 19'b0100010000000000_100;
      patterns[1300] = 19'b1000010000000100_100;
      patterns[1301] = 19'b1001010000000100_100;
      patterns[1302] = 19'b1010010000000100_100;
      patterns[1303] = 19'b1011010000000100_100;
      patterns[1304] = 19'b0100010000000000_100;
      patterns[1305] = 19'b1000010000000101_101;
      patterns[1306] = 19'b1001010000000101_101;
      patterns[1307] = 19'b1010010000000101_101;
      patterns[1308] = 19'b1011010000000101_101;
      patterns[1309] = 19'b0100010000000000_100;
      patterns[1310] = 19'b1000010000000110_110;
      patterns[1311] = 19'b1001010000000110_110;
      patterns[1312] = 19'b1010010000000110_110;
      patterns[1313] = 19'b1011010000000110_110;
      patterns[1314] = 19'b0100010000000000_100;
      patterns[1315] = 19'b1000010000000111_111;
      patterns[1316] = 19'b1001010000000111_111;
      patterns[1317] = 19'b1010010000000111_111;
      patterns[1318] = 19'b1011010000000111_111;
      patterns[1319] = 19'b0100010000000000_100;
      patterns[1320] = 19'b1000010000010000_000;
      patterns[1321] = 19'b1001010000010000_000;
      patterns[1322] = 19'b1010010000010000_000;
      patterns[1323] = 19'b1011010000010000_000;
      patterns[1324] = 19'b0100010000010000_100;
      patterns[1325] = 19'b1000010000010001_001;
      patterns[1326] = 19'b1001010000010001_001;
      patterns[1327] = 19'b1010010000010001_001;
      patterns[1328] = 19'b1011010000010001_001;
      patterns[1329] = 19'b0100010000010000_100;
      patterns[1330] = 19'b1000010000010010_010;
      patterns[1331] = 19'b1001010000010010_010;
      patterns[1332] = 19'b1010010000010010_010;
      patterns[1333] = 19'b1011010000010010_010;
      patterns[1334] = 19'b0100010000010000_100;
      patterns[1335] = 19'b1000010000010011_011;
      patterns[1336] = 19'b1001010000010011_011;
      patterns[1337] = 19'b1010010000010011_011;
      patterns[1338] = 19'b1011010000010011_011;
      patterns[1339] = 19'b0100010000010000_100;
      patterns[1340] = 19'b1000010000010100_100;
      patterns[1341] = 19'b1001010000010100_100;
      patterns[1342] = 19'b1010010000010100_100;
      patterns[1343] = 19'b1011010000010100_100;
      patterns[1344] = 19'b0100010000010000_100;
      patterns[1345] = 19'b1000010000010101_101;
      patterns[1346] = 19'b1001010000010101_101;
      patterns[1347] = 19'b1010010000010101_101;
      patterns[1348] = 19'b1011010000010101_101;
      patterns[1349] = 19'b0100010000010000_100;
      patterns[1350] = 19'b1000010000010110_110;
      patterns[1351] = 19'b1001010000010110_110;
      patterns[1352] = 19'b1010010000010110_110;
      patterns[1353] = 19'b1011010000010110_110;
      patterns[1354] = 19'b0100010000010000_100;
      patterns[1355] = 19'b1000010000010111_111;
      patterns[1356] = 19'b1001010000010111_111;
      patterns[1357] = 19'b1010010000010111_111;
      patterns[1358] = 19'b1011010000010111_111;
      patterns[1359] = 19'b0100010000010000_100;
      patterns[1360] = 19'b1000010000100000_000;
      patterns[1361] = 19'b1001010000100000_000;
      patterns[1362] = 19'b1010010000100000_000;
      patterns[1363] = 19'b1011010000100000_000;
      patterns[1364] = 19'b0100010000100000_100;
      patterns[1365] = 19'b1000010000100001_001;
      patterns[1366] = 19'b1001010000100001_001;
      patterns[1367] = 19'b1010010000100001_001;
      patterns[1368] = 19'b1011010000100001_001;
      patterns[1369] = 19'b0100010000100000_100;
      patterns[1370] = 19'b1000010000100010_010;
      patterns[1371] = 19'b1001010000100010_010;
      patterns[1372] = 19'b1010010000100010_010;
      patterns[1373] = 19'b1011010000100010_010;
      patterns[1374] = 19'b0100010000100000_100;
      patterns[1375] = 19'b1000010000100011_011;
      patterns[1376] = 19'b1001010000100011_011;
      patterns[1377] = 19'b1010010000100011_011;
      patterns[1378] = 19'b1011010000100011_011;
      patterns[1379] = 19'b0100010000100000_100;
      patterns[1380] = 19'b1000010000100100_100;
      patterns[1381] = 19'b1001010000100100_100;
      patterns[1382] = 19'b1010010000100100_100;
      patterns[1383] = 19'b1011010000100100_100;
      patterns[1384] = 19'b0100010000100000_100;
      patterns[1385] = 19'b1000010000100101_101;
      patterns[1386] = 19'b1001010000100101_101;
      patterns[1387] = 19'b1010010000100101_101;
      patterns[1388] = 19'b1011010000100101_101;
      patterns[1389] = 19'b0100010000100000_100;
      patterns[1390] = 19'b1000010000100110_110;
      patterns[1391] = 19'b1001010000100110_110;
      patterns[1392] = 19'b1010010000100110_110;
      patterns[1393] = 19'b1011010000100110_110;
      patterns[1394] = 19'b0100010000100000_100;
      patterns[1395] = 19'b1000010000100111_111;
      patterns[1396] = 19'b1001010000100111_111;
      patterns[1397] = 19'b1010010000100111_111;
      patterns[1398] = 19'b1011010000100111_111;
      patterns[1399] = 19'b0100010000100000_100;
      patterns[1400] = 19'b1000010000110000_000;
      patterns[1401] = 19'b1001010000110000_000;
      patterns[1402] = 19'b1010010000110000_000;
      patterns[1403] = 19'b1011010000110000_000;
      patterns[1404] = 19'b0100010000110000_100;
      patterns[1405] = 19'b1000010000110001_001;
      patterns[1406] = 19'b1001010000110001_001;
      patterns[1407] = 19'b1010010000110001_001;
      patterns[1408] = 19'b1011010000110001_001;
      patterns[1409] = 19'b0100010000110000_100;
      patterns[1410] = 19'b1000010000110010_010;
      patterns[1411] = 19'b1001010000110010_010;
      patterns[1412] = 19'b1010010000110010_010;
      patterns[1413] = 19'b1011010000110010_010;
      patterns[1414] = 19'b0100010000110000_100;
      patterns[1415] = 19'b1000010000110011_011;
      patterns[1416] = 19'b1001010000110011_011;
      patterns[1417] = 19'b1010010000110011_011;
      patterns[1418] = 19'b1011010000110011_011;
      patterns[1419] = 19'b0100010000110000_100;
      patterns[1420] = 19'b1000010000110100_100;
      patterns[1421] = 19'b1001010000110100_100;
      patterns[1422] = 19'b1010010000110100_100;
      patterns[1423] = 19'b1011010000110100_100;
      patterns[1424] = 19'b0100010000110000_100;
      patterns[1425] = 19'b1000010000110101_101;
      patterns[1426] = 19'b1001010000110101_101;
      patterns[1427] = 19'b1010010000110101_101;
      patterns[1428] = 19'b1011010000110101_101;
      patterns[1429] = 19'b0100010000110000_100;
      patterns[1430] = 19'b1000010000110110_110;
      patterns[1431] = 19'b1001010000110110_110;
      patterns[1432] = 19'b1010010000110110_110;
      patterns[1433] = 19'b1011010000110110_110;
      patterns[1434] = 19'b0100010000110000_100;
      patterns[1435] = 19'b1000010000110111_111;
      patterns[1436] = 19'b1001010000110111_111;
      patterns[1437] = 19'b1010010000110111_111;
      patterns[1438] = 19'b1011010000110111_111;
      patterns[1439] = 19'b0100010000110000_100;
      patterns[1440] = 19'b1000010001000000_000;
      patterns[1441] = 19'b1001010001000000_000;
      patterns[1442] = 19'b1010010001000000_000;
      patterns[1443] = 19'b1011010001000000_000;
      patterns[1444] = 19'b0100010001000000_100;
      patterns[1445] = 19'b1000010001000001_001;
      patterns[1446] = 19'b1001010001000001_001;
      patterns[1447] = 19'b1010010001000001_001;
      patterns[1448] = 19'b1011010001000001_001;
      patterns[1449] = 19'b0100010001000000_100;
      patterns[1450] = 19'b1000010001000010_010;
      patterns[1451] = 19'b1001010001000010_010;
      patterns[1452] = 19'b1010010001000010_010;
      patterns[1453] = 19'b1011010001000010_010;
      patterns[1454] = 19'b0100010001000000_100;
      patterns[1455] = 19'b1000010001000011_011;
      patterns[1456] = 19'b1001010001000011_011;
      patterns[1457] = 19'b1010010001000011_011;
      patterns[1458] = 19'b1011010001000011_011;
      patterns[1459] = 19'b0100010001000000_100;
      patterns[1460] = 19'b1000010001000100_100;
      patterns[1461] = 19'b1001010001000100_100;
      patterns[1462] = 19'b1010010001000100_100;
      patterns[1463] = 19'b1011010001000100_100;
      patterns[1464] = 19'b0100010001000000_100;
      patterns[1465] = 19'b1000010001000101_101;
      patterns[1466] = 19'b1001010001000101_101;
      patterns[1467] = 19'b1010010001000101_101;
      patterns[1468] = 19'b1011010001000101_101;
      patterns[1469] = 19'b0100010001000000_100;
      patterns[1470] = 19'b1000010001000110_110;
      patterns[1471] = 19'b1001010001000110_110;
      patterns[1472] = 19'b1010010001000110_110;
      patterns[1473] = 19'b1011010001000110_110;
      patterns[1474] = 19'b0100010001000000_100;
      patterns[1475] = 19'b1000010001000111_111;
      patterns[1476] = 19'b1001010001000111_111;
      patterns[1477] = 19'b1010010001000111_111;
      patterns[1478] = 19'b1011010001000111_111;
      patterns[1479] = 19'b0100010001000000_100;
      patterns[1480] = 19'b1000010001010000_000;
      patterns[1481] = 19'b1001010001010000_000;
      patterns[1482] = 19'b1010010001010000_000;
      patterns[1483] = 19'b1011010001010000_000;
      patterns[1484] = 19'b0100010001010000_100;
      patterns[1485] = 19'b1000010001010001_001;
      patterns[1486] = 19'b1001010001010001_001;
      patterns[1487] = 19'b1010010001010001_001;
      patterns[1488] = 19'b1011010001010001_001;
      patterns[1489] = 19'b0100010001010000_100;
      patterns[1490] = 19'b1000010001010010_010;
      patterns[1491] = 19'b1001010001010010_010;
      patterns[1492] = 19'b1010010001010010_010;
      patterns[1493] = 19'b1011010001010010_010;
      patterns[1494] = 19'b0100010001010000_100;
      patterns[1495] = 19'b1000010001010011_011;
      patterns[1496] = 19'b1001010001010011_011;
      patterns[1497] = 19'b1010010001010011_011;
      patterns[1498] = 19'b1011010001010011_011;
      patterns[1499] = 19'b0100010001010000_100;
      patterns[1500] = 19'b1000010001010100_100;
      patterns[1501] = 19'b1001010001010100_100;
      patterns[1502] = 19'b1010010001010100_100;
      patterns[1503] = 19'b1011010001010100_100;
      patterns[1504] = 19'b0100010001010000_100;
      patterns[1505] = 19'b1000010001010101_101;
      patterns[1506] = 19'b1001010001010101_101;
      patterns[1507] = 19'b1010010001010101_101;
      patterns[1508] = 19'b1011010001010101_101;
      patterns[1509] = 19'b0100010001010000_100;
      patterns[1510] = 19'b1000010001010110_110;
      patterns[1511] = 19'b1001010001010110_110;
      patterns[1512] = 19'b1010010001010110_110;
      patterns[1513] = 19'b1011010001010110_110;
      patterns[1514] = 19'b0100010001010000_100;
      patterns[1515] = 19'b1000010001010111_111;
      patterns[1516] = 19'b1001010001010111_111;
      patterns[1517] = 19'b1010010001010111_111;
      patterns[1518] = 19'b1011010001010111_111;
      patterns[1519] = 19'b0100010001010000_100;
      patterns[1520] = 19'b1000010001100000_000;
      patterns[1521] = 19'b1001010001100000_000;
      patterns[1522] = 19'b1010010001100000_000;
      patterns[1523] = 19'b1011010001100000_000;
      patterns[1524] = 19'b0100010001100000_100;
      patterns[1525] = 19'b1000010001100001_001;
      patterns[1526] = 19'b1001010001100001_001;
      patterns[1527] = 19'b1010010001100001_001;
      patterns[1528] = 19'b1011010001100001_001;
      patterns[1529] = 19'b0100010001100000_100;
      patterns[1530] = 19'b1000010001100010_010;
      patterns[1531] = 19'b1001010001100010_010;
      patterns[1532] = 19'b1010010001100010_010;
      patterns[1533] = 19'b1011010001100010_010;
      patterns[1534] = 19'b0100010001100000_100;
      patterns[1535] = 19'b1000010001100011_011;
      patterns[1536] = 19'b1001010001100011_011;
      patterns[1537] = 19'b1010010001100011_011;
      patterns[1538] = 19'b1011010001100011_011;
      patterns[1539] = 19'b0100010001100000_100;
      patterns[1540] = 19'b1000010001100100_100;
      patterns[1541] = 19'b1001010001100100_100;
      patterns[1542] = 19'b1010010001100100_100;
      patterns[1543] = 19'b1011010001100100_100;
      patterns[1544] = 19'b0100010001100000_100;
      patterns[1545] = 19'b1000010001100101_101;
      patterns[1546] = 19'b1001010001100101_101;
      patterns[1547] = 19'b1010010001100101_101;
      patterns[1548] = 19'b1011010001100101_101;
      patterns[1549] = 19'b0100010001100000_100;
      patterns[1550] = 19'b1000010001100110_110;
      patterns[1551] = 19'b1001010001100110_110;
      patterns[1552] = 19'b1010010001100110_110;
      patterns[1553] = 19'b1011010001100110_110;
      patterns[1554] = 19'b0100010001100000_100;
      patterns[1555] = 19'b1000010001100111_111;
      patterns[1556] = 19'b1001010001100111_111;
      patterns[1557] = 19'b1010010001100111_111;
      patterns[1558] = 19'b1011010001100111_111;
      patterns[1559] = 19'b0100010001100000_100;
      patterns[1560] = 19'b1000010001110000_000;
      patterns[1561] = 19'b1001010001110000_000;
      patterns[1562] = 19'b1010010001110000_000;
      patterns[1563] = 19'b1011010001110000_000;
      patterns[1564] = 19'b0100010001110000_100;
      patterns[1565] = 19'b1000010001110001_001;
      patterns[1566] = 19'b1001010001110001_001;
      patterns[1567] = 19'b1010010001110001_001;
      patterns[1568] = 19'b1011010001110001_001;
      patterns[1569] = 19'b0100010001110000_100;
      patterns[1570] = 19'b1000010001110010_010;
      patterns[1571] = 19'b1001010001110010_010;
      patterns[1572] = 19'b1010010001110010_010;
      patterns[1573] = 19'b1011010001110010_010;
      patterns[1574] = 19'b0100010001110000_100;
      patterns[1575] = 19'b1000010001110011_011;
      patterns[1576] = 19'b1001010001110011_011;
      patterns[1577] = 19'b1010010001110011_011;
      patterns[1578] = 19'b1011010001110011_011;
      patterns[1579] = 19'b0100010001110000_100;
      patterns[1580] = 19'b1000010001110100_100;
      patterns[1581] = 19'b1001010001110100_100;
      patterns[1582] = 19'b1010010001110100_100;
      patterns[1583] = 19'b1011010001110100_100;
      patterns[1584] = 19'b0100010001110000_100;
      patterns[1585] = 19'b1000010001110101_101;
      patterns[1586] = 19'b1001010001110101_101;
      patterns[1587] = 19'b1010010001110101_101;
      patterns[1588] = 19'b1011010001110101_101;
      patterns[1589] = 19'b0100010001110000_100;
      patterns[1590] = 19'b1000010001110110_110;
      patterns[1591] = 19'b1001010001110110_110;
      patterns[1592] = 19'b1010010001110110_110;
      patterns[1593] = 19'b1011010001110110_110;
      patterns[1594] = 19'b0100010001110000_100;
      patterns[1595] = 19'b1000010001110111_111;
      patterns[1596] = 19'b1001010001110111_111;
      patterns[1597] = 19'b1010010001110111_111;
      patterns[1598] = 19'b1011010001110111_111;
      patterns[1599] = 19'b0100010001110000_100;
      patterns[1600] = 19'b1000010100000000_000;
      patterns[1601] = 19'b1001010100000000_000;
      patterns[1602] = 19'b1010010100000000_000;
      patterns[1603] = 19'b1011010100000000_000;
      patterns[1604] = 19'b0100010100000000_101;
      patterns[1605] = 19'b1000010100000001_001;
      patterns[1606] = 19'b1001010100000001_001;
      patterns[1607] = 19'b1010010100000001_001;
      patterns[1608] = 19'b1011010100000001_001;
      patterns[1609] = 19'b0100010100000000_101;
      patterns[1610] = 19'b1000010100000010_010;
      patterns[1611] = 19'b1001010100000010_010;
      patterns[1612] = 19'b1010010100000010_010;
      patterns[1613] = 19'b1011010100000010_010;
      patterns[1614] = 19'b0100010100000000_101;
      patterns[1615] = 19'b1000010100000011_011;
      patterns[1616] = 19'b1001010100000011_011;
      patterns[1617] = 19'b1010010100000011_011;
      patterns[1618] = 19'b1011010100000011_011;
      patterns[1619] = 19'b0100010100000000_101;
      patterns[1620] = 19'b1000010100000100_100;
      patterns[1621] = 19'b1001010100000100_100;
      patterns[1622] = 19'b1010010100000100_100;
      patterns[1623] = 19'b1011010100000100_100;
      patterns[1624] = 19'b0100010100000000_101;
      patterns[1625] = 19'b1000010100000101_101;
      patterns[1626] = 19'b1001010100000101_101;
      patterns[1627] = 19'b1010010100000101_101;
      patterns[1628] = 19'b1011010100000101_101;
      patterns[1629] = 19'b0100010100000000_101;
      patterns[1630] = 19'b1000010100000110_110;
      patterns[1631] = 19'b1001010100000110_110;
      patterns[1632] = 19'b1010010100000110_110;
      patterns[1633] = 19'b1011010100000110_110;
      patterns[1634] = 19'b0100010100000000_101;
      patterns[1635] = 19'b1000010100000111_111;
      patterns[1636] = 19'b1001010100000111_111;
      patterns[1637] = 19'b1010010100000111_111;
      patterns[1638] = 19'b1011010100000111_111;
      patterns[1639] = 19'b0100010100000000_101;
      patterns[1640] = 19'b1000010100010000_000;
      patterns[1641] = 19'b1001010100010000_000;
      patterns[1642] = 19'b1010010100010000_000;
      patterns[1643] = 19'b1011010100010000_000;
      patterns[1644] = 19'b0100010100010000_101;
      patterns[1645] = 19'b1000010100010001_001;
      patterns[1646] = 19'b1001010100010001_001;
      patterns[1647] = 19'b1010010100010001_001;
      patterns[1648] = 19'b1011010100010001_001;
      patterns[1649] = 19'b0100010100010000_101;
      patterns[1650] = 19'b1000010100010010_010;
      patterns[1651] = 19'b1001010100010010_010;
      patterns[1652] = 19'b1010010100010010_010;
      patterns[1653] = 19'b1011010100010010_010;
      patterns[1654] = 19'b0100010100010000_101;
      patterns[1655] = 19'b1000010100010011_011;
      patterns[1656] = 19'b1001010100010011_011;
      patterns[1657] = 19'b1010010100010011_011;
      patterns[1658] = 19'b1011010100010011_011;
      patterns[1659] = 19'b0100010100010000_101;
      patterns[1660] = 19'b1000010100010100_100;
      patterns[1661] = 19'b1001010100010100_100;
      patterns[1662] = 19'b1010010100010100_100;
      patterns[1663] = 19'b1011010100010100_100;
      patterns[1664] = 19'b0100010100010000_101;
      patterns[1665] = 19'b1000010100010101_101;
      patterns[1666] = 19'b1001010100010101_101;
      patterns[1667] = 19'b1010010100010101_101;
      patterns[1668] = 19'b1011010100010101_101;
      patterns[1669] = 19'b0100010100010000_101;
      patterns[1670] = 19'b1000010100010110_110;
      patterns[1671] = 19'b1001010100010110_110;
      patterns[1672] = 19'b1010010100010110_110;
      patterns[1673] = 19'b1011010100010110_110;
      patterns[1674] = 19'b0100010100010000_101;
      patterns[1675] = 19'b1000010100010111_111;
      patterns[1676] = 19'b1001010100010111_111;
      patterns[1677] = 19'b1010010100010111_111;
      patterns[1678] = 19'b1011010100010111_111;
      patterns[1679] = 19'b0100010100010000_101;
      patterns[1680] = 19'b1000010100100000_000;
      patterns[1681] = 19'b1001010100100000_000;
      patterns[1682] = 19'b1010010100100000_000;
      patterns[1683] = 19'b1011010100100000_000;
      patterns[1684] = 19'b0100010100100000_101;
      patterns[1685] = 19'b1000010100100001_001;
      patterns[1686] = 19'b1001010100100001_001;
      patterns[1687] = 19'b1010010100100001_001;
      patterns[1688] = 19'b1011010100100001_001;
      patterns[1689] = 19'b0100010100100000_101;
      patterns[1690] = 19'b1000010100100010_010;
      patterns[1691] = 19'b1001010100100010_010;
      patterns[1692] = 19'b1010010100100010_010;
      patterns[1693] = 19'b1011010100100010_010;
      patterns[1694] = 19'b0100010100100000_101;
      patterns[1695] = 19'b1000010100100011_011;
      patterns[1696] = 19'b1001010100100011_011;
      patterns[1697] = 19'b1010010100100011_011;
      patterns[1698] = 19'b1011010100100011_011;
      patterns[1699] = 19'b0100010100100000_101;
      patterns[1700] = 19'b1000010100100100_100;
      patterns[1701] = 19'b1001010100100100_100;
      patterns[1702] = 19'b1010010100100100_100;
      patterns[1703] = 19'b1011010100100100_100;
      patterns[1704] = 19'b0100010100100000_101;
      patterns[1705] = 19'b1000010100100101_101;
      patterns[1706] = 19'b1001010100100101_101;
      patterns[1707] = 19'b1010010100100101_101;
      patterns[1708] = 19'b1011010100100101_101;
      patterns[1709] = 19'b0100010100100000_101;
      patterns[1710] = 19'b1000010100100110_110;
      patterns[1711] = 19'b1001010100100110_110;
      patterns[1712] = 19'b1010010100100110_110;
      patterns[1713] = 19'b1011010100100110_110;
      patterns[1714] = 19'b0100010100100000_101;
      patterns[1715] = 19'b1000010100100111_111;
      patterns[1716] = 19'b1001010100100111_111;
      patterns[1717] = 19'b1010010100100111_111;
      patterns[1718] = 19'b1011010100100111_111;
      patterns[1719] = 19'b0100010100100000_101;
      patterns[1720] = 19'b1000010100110000_000;
      patterns[1721] = 19'b1001010100110000_000;
      patterns[1722] = 19'b1010010100110000_000;
      patterns[1723] = 19'b1011010100110000_000;
      patterns[1724] = 19'b0100010100110000_101;
      patterns[1725] = 19'b1000010100110001_001;
      patterns[1726] = 19'b1001010100110001_001;
      patterns[1727] = 19'b1010010100110001_001;
      patterns[1728] = 19'b1011010100110001_001;
      patterns[1729] = 19'b0100010100110000_101;
      patterns[1730] = 19'b1000010100110010_010;
      patterns[1731] = 19'b1001010100110010_010;
      patterns[1732] = 19'b1010010100110010_010;
      patterns[1733] = 19'b1011010100110010_010;
      patterns[1734] = 19'b0100010100110000_101;
      patterns[1735] = 19'b1000010100110011_011;
      patterns[1736] = 19'b1001010100110011_011;
      patterns[1737] = 19'b1010010100110011_011;
      patterns[1738] = 19'b1011010100110011_011;
      patterns[1739] = 19'b0100010100110000_101;
      patterns[1740] = 19'b1000010100110100_100;
      patterns[1741] = 19'b1001010100110100_100;
      patterns[1742] = 19'b1010010100110100_100;
      patterns[1743] = 19'b1011010100110100_100;
      patterns[1744] = 19'b0100010100110000_101;
      patterns[1745] = 19'b1000010100110101_101;
      patterns[1746] = 19'b1001010100110101_101;
      patterns[1747] = 19'b1010010100110101_101;
      patterns[1748] = 19'b1011010100110101_101;
      patterns[1749] = 19'b0100010100110000_101;
      patterns[1750] = 19'b1000010100110110_110;
      patterns[1751] = 19'b1001010100110110_110;
      patterns[1752] = 19'b1010010100110110_110;
      patterns[1753] = 19'b1011010100110110_110;
      patterns[1754] = 19'b0100010100110000_101;
      patterns[1755] = 19'b1000010100110111_111;
      patterns[1756] = 19'b1001010100110111_111;
      patterns[1757] = 19'b1010010100110111_111;
      patterns[1758] = 19'b1011010100110111_111;
      patterns[1759] = 19'b0100010100110000_101;
      patterns[1760] = 19'b1000010101000000_000;
      patterns[1761] = 19'b1001010101000000_000;
      patterns[1762] = 19'b1010010101000000_000;
      patterns[1763] = 19'b1011010101000000_000;
      patterns[1764] = 19'b0100010101000000_101;
      patterns[1765] = 19'b1000010101000001_001;
      patterns[1766] = 19'b1001010101000001_001;
      patterns[1767] = 19'b1010010101000001_001;
      patterns[1768] = 19'b1011010101000001_001;
      patterns[1769] = 19'b0100010101000000_101;
      patterns[1770] = 19'b1000010101000010_010;
      patterns[1771] = 19'b1001010101000010_010;
      patterns[1772] = 19'b1010010101000010_010;
      patterns[1773] = 19'b1011010101000010_010;
      patterns[1774] = 19'b0100010101000000_101;
      patterns[1775] = 19'b1000010101000011_011;
      patterns[1776] = 19'b1001010101000011_011;
      patterns[1777] = 19'b1010010101000011_011;
      patterns[1778] = 19'b1011010101000011_011;
      patterns[1779] = 19'b0100010101000000_101;
      patterns[1780] = 19'b1000010101000100_100;
      patterns[1781] = 19'b1001010101000100_100;
      patterns[1782] = 19'b1010010101000100_100;
      patterns[1783] = 19'b1011010101000100_100;
      patterns[1784] = 19'b0100010101000000_101;
      patterns[1785] = 19'b1000010101000101_101;
      patterns[1786] = 19'b1001010101000101_101;
      patterns[1787] = 19'b1010010101000101_101;
      patterns[1788] = 19'b1011010101000101_101;
      patterns[1789] = 19'b0100010101000000_101;
      patterns[1790] = 19'b1000010101000110_110;
      patterns[1791] = 19'b1001010101000110_110;
      patterns[1792] = 19'b1010010101000110_110;
      patterns[1793] = 19'b1011010101000110_110;
      patterns[1794] = 19'b0100010101000000_101;
      patterns[1795] = 19'b1000010101000111_111;
      patterns[1796] = 19'b1001010101000111_111;
      patterns[1797] = 19'b1010010101000111_111;
      patterns[1798] = 19'b1011010101000111_111;
      patterns[1799] = 19'b0100010101000000_101;
      patterns[1800] = 19'b1000010101010000_000;
      patterns[1801] = 19'b1001010101010000_000;
      patterns[1802] = 19'b1010010101010000_000;
      patterns[1803] = 19'b1011010101010000_000;
      patterns[1804] = 19'b0100010101010000_101;
      patterns[1805] = 19'b1000010101010001_001;
      patterns[1806] = 19'b1001010101010001_001;
      patterns[1807] = 19'b1010010101010001_001;
      patterns[1808] = 19'b1011010101010001_001;
      patterns[1809] = 19'b0100010101010000_101;
      patterns[1810] = 19'b1000010101010010_010;
      patterns[1811] = 19'b1001010101010010_010;
      patterns[1812] = 19'b1010010101010010_010;
      patterns[1813] = 19'b1011010101010010_010;
      patterns[1814] = 19'b0100010101010000_101;
      patterns[1815] = 19'b1000010101010011_011;
      patterns[1816] = 19'b1001010101010011_011;
      patterns[1817] = 19'b1010010101010011_011;
      patterns[1818] = 19'b1011010101010011_011;
      patterns[1819] = 19'b0100010101010000_101;
      patterns[1820] = 19'b1000010101010100_100;
      patterns[1821] = 19'b1001010101010100_100;
      patterns[1822] = 19'b1010010101010100_100;
      patterns[1823] = 19'b1011010101010100_100;
      patterns[1824] = 19'b0100010101010000_101;
      patterns[1825] = 19'b1000010101010101_101;
      patterns[1826] = 19'b1001010101010101_101;
      patterns[1827] = 19'b1010010101010101_101;
      patterns[1828] = 19'b1011010101010101_101;
      patterns[1829] = 19'b0100010101010000_101;
      patterns[1830] = 19'b1000010101010110_110;
      patterns[1831] = 19'b1001010101010110_110;
      patterns[1832] = 19'b1010010101010110_110;
      patterns[1833] = 19'b1011010101010110_110;
      patterns[1834] = 19'b0100010101010000_101;
      patterns[1835] = 19'b1000010101010111_111;
      patterns[1836] = 19'b1001010101010111_111;
      patterns[1837] = 19'b1010010101010111_111;
      patterns[1838] = 19'b1011010101010111_111;
      patterns[1839] = 19'b0100010101010000_101;
      patterns[1840] = 19'b1000010101100000_000;
      patterns[1841] = 19'b1001010101100000_000;
      patterns[1842] = 19'b1010010101100000_000;
      patterns[1843] = 19'b1011010101100000_000;
      patterns[1844] = 19'b0100010101100000_101;
      patterns[1845] = 19'b1000010101100001_001;
      patterns[1846] = 19'b1001010101100001_001;
      patterns[1847] = 19'b1010010101100001_001;
      patterns[1848] = 19'b1011010101100001_001;
      patterns[1849] = 19'b0100010101100000_101;
      patterns[1850] = 19'b1000010101100010_010;
      patterns[1851] = 19'b1001010101100010_010;
      patterns[1852] = 19'b1010010101100010_010;
      patterns[1853] = 19'b1011010101100010_010;
      patterns[1854] = 19'b0100010101100000_101;
      patterns[1855] = 19'b1000010101100011_011;
      patterns[1856] = 19'b1001010101100011_011;
      patterns[1857] = 19'b1010010101100011_011;
      patterns[1858] = 19'b1011010101100011_011;
      patterns[1859] = 19'b0100010101100000_101;
      patterns[1860] = 19'b1000010101100100_100;
      patterns[1861] = 19'b1001010101100100_100;
      patterns[1862] = 19'b1010010101100100_100;
      patterns[1863] = 19'b1011010101100100_100;
      patterns[1864] = 19'b0100010101100000_101;
      patterns[1865] = 19'b1000010101100101_101;
      patterns[1866] = 19'b1001010101100101_101;
      patterns[1867] = 19'b1010010101100101_101;
      patterns[1868] = 19'b1011010101100101_101;
      patterns[1869] = 19'b0100010101100000_101;
      patterns[1870] = 19'b1000010101100110_110;
      patterns[1871] = 19'b1001010101100110_110;
      patterns[1872] = 19'b1010010101100110_110;
      patterns[1873] = 19'b1011010101100110_110;
      patterns[1874] = 19'b0100010101100000_101;
      patterns[1875] = 19'b1000010101100111_111;
      patterns[1876] = 19'b1001010101100111_111;
      patterns[1877] = 19'b1010010101100111_111;
      patterns[1878] = 19'b1011010101100111_111;
      patterns[1879] = 19'b0100010101100000_101;
      patterns[1880] = 19'b1000010101110000_000;
      patterns[1881] = 19'b1001010101110000_000;
      patterns[1882] = 19'b1010010101110000_000;
      patterns[1883] = 19'b1011010101110000_000;
      patterns[1884] = 19'b0100010101110000_101;
      patterns[1885] = 19'b1000010101110001_001;
      patterns[1886] = 19'b1001010101110001_001;
      patterns[1887] = 19'b1010010101110001_001;
      patterns[1888] = 19'b1011010101110001_001;
      patterns[1889] = 19'b0100010101110000_101;
      patterns[1890] = 19'b1000010101110010_010;
      patterns[1891] = 19'b1001010101110010_010;
      patterns[1892] = 19'b1010010101110010_010;
      patterns[1893] = 19'b1011010101110010_010;
      patterns[1894] = 19'b0100010101110000_101;
      patterns[1895] = 19'b1000010101110011_011;
      patterns[1896] = 19'b1001010101110011_011;
      patterns[1897] = 19'b1010010101110011_011;
      patterns[1898] = 19'b1011010101110011_011;
      patterns[1899] = 19'b0100010101110000_101;
      patterns[1900] = 19'b1000010101110100_100;
      patterns[1901] = 19'b1001010101110100_100;
      patterns[1902] = 19'b1010010101110100_100;
      patterns[1903] = 19'b1011010101110100_100;
      patterns[1904] = 19'b0100010101110000_101;
      patterns[1905] = 19'b1000010101110101_101;
      patterns[1906] = 19'b1001010101110101_101;
      patterns[1907] = 19'b1010010101110101_101;
      patterns[1908] = 19'b1011010101110101_101;
      patterns[1909] = 19'b0100010101110000_101;
      patterns[1910] = 19'b1000010101110110_110;
      patterns[1911] = 19'b1001010101110110_110;
      patterns[1912] = 19'b1010010101110110_110;
      patterns[1913] = 19'b1011010101110110_110;
      patterns[1914] = 19'b0100010101110000_101;
      patterns[1915] = 19'b1000010101110111_111;
      patterns[1916] = 19'b1001010101110111_111;
      patterns[1917] = 19'b1010010101110111_111;
      patterns[1918] = 19'b1011010101110111_111;
      patterns[1919] = 19'b0100010101110000_101;
      patterns[1920] = 19'b1000011000000000_000;
      patterns[1921] = 19'b1001011000000000_000;
      patterns[1922] = 19'b1010011000000000_000;
      patterns[1923] = 19'b1011011000000000_000;
      patterns[1924] = 19'b0100011000000000_110;
      patterns[1925] = 19'b1000011000000001_001;
      patterns[1926] = 19'b1001011000000001_001;
      patterns[1927] = 19'b1010011000000001_001;
      patterns[1928] = 19'b1011011000000001_001;
      patterns[1929] = 19'b0100011000000000_110;
      patterns[1930] = 19'b1000011000000010_010;
      patterns[1931] = 19'b1001011000000010_010;
      patterns[1932] = 19'b1010011000000010_010;
      patterns[1933] = 19'b1011011000000010_010;
      patterns[1934] = 19'b0100011000000000_110;
      patterns[1935] = 19'b1000011000000011_011;
      patterns[1936] = 19'b1001011000000011_011;
      patterns[1937] = 19'b1010011000000011_011;
      patterns[1938] = 19'b1011011000000011_011;
      patterns[1939] = 19'b0100011000000000_110;
      patterns[1940] = 19'b1000011000000100_100;
      patterns[1941] = 19'b1001011000000100_100;
      patterns[1942] = 19'b1010011000000100_100;
      patterns[1943] = 19'b1011011000000100_100;
      patterns[1944] = 19'b0100011000000000_110;
      patterns[1945] = 19'b1000011000000101_101;
      patterns[1946] = 19'b1001011000000101_101;
      patterns[1947] = 19'b1010011000000101_101;
      patterns[1948] = 19'b1011011000000101_101;
      patterns[1949] = 19'b0100011000000000_110;
      patterns[1950] = 19'b1000011000000110_110;
      patterns[1951] = 19'b1001011000000110_110;
      patterns[1952] = 19'b1010011000000110_110;
      patterns[1953] = 19'b1011011000000110_110;
      patterns[1954] = 19'b0100011000000000_110;
      patterns[1955] = 19'b1000011000000111_111;
      patterns[1956] = 19'b1001011000000111_111;
      patterns[1957] = 19'b1010011000000111_111;
      patterns[1958] = 19'b1011011000000111_111;
      patterns[1959] = 19'b0100011000000000_110;
      patterns[1960] = 19'b1000011000010000_000;
      patterns[1961] = 19'b1001011000010000_000;
      patterns[1962] = 19'b1010011000010000_000;
      patterns[1963] = 19'b1011011000010000_000;
      patterns[1964] = 19'b0100011000010000_110;
      patterns[1965] = 19'b1000011000010001_001;
      patterns[1966] = 19'b1001011000010001_001;
      patterns[1967] = 19'b1010011000010001_001;
      patterns[1968] = 19'b1011011000010001_001;
      patterns[1969] = 19'b0100011000010000_110;
      patterns[1970] = 19'b1000011000010010_010;
      patterns[1971] = 19'b1001011000010010_010;
      patterns[1972] = 19'b1010011000010010_010;
      patterns[1973] = 19'b1011011000010010_010;
      patterns[1974] = 19'b0100011000010000_110;
      patterns[1975] = 19'b1000011000010011_011;
      patterns[1976] = 19'b1001011000010011_011;
      patterns[1977] = 19'b1010011000010011_011;
      patterns[1978] = 19'b1011011000010011_011;
      patterns[1979] = 19'b0100011000010000_110;
      patterns[1980] = 19'b1000011000010100_100;
      patterns[1981] = 19'b1001011000010100_100;
      patterns[1982] = 19'b1010011000010100_100;
      patterns[1983] = 19'b1011011000010100_100;
      patterns[1984] = 19'b0100011000010000_110;
      patterns[1985] = 19'b1000011000010101_101;
      patterns[1986] = 19'b1001011000010101_101;
      patterns[1987] = 19'b1010011000010101_101;
      patterns[1988] = 19'b1011011000010101_101;
      patterns[1989] = 19'b0100011000010000_110;
      patterns[1990] = 19'b1000011000010110_110;
      patterns[1991] = 19'b1001011000010110_110;
      patterns[1992] = 19'b1010011000010110_110;
      patterns[1993] = 19'b1011011000010110_110;
      patterns[1994] = 19'b0100011000010000_110;
      patterns[1995] = 19'b1000011000010111_111;
      patterns[1996] = 19'b1001011000010111_111;
      patterns[1997] = 19'b1010011000010111_111;
      patterns[1998] = 19'b1011011000010111_111;
      patterns[1999] = 19'b0100011000010000_110;
      patterns[2000] = 19'b1000011000100000_000;
      patterns[2001] = 19'b1001011000100000_000;
      patterns[2002] = 19'b1010011000100000_000;
      patterns[2003] = 19'b1011011000100000_000;
      patterns[2004] = 19'b0100011000100000_110;
      patterns[2005] = 19'b1000011000100001_001;
      patterns[2006] = 19'b1001011000100001_001;
      patterns[2007] = 19'b1010011000100001_001;
      patterns[2008] = 19'b1011011000100001_001;
      patterns[2009] = 19'b0100011000100000_110;
      patterns[2010] = 19'b1000011000100010_010;
      patterns[2011] = 19'b1001011000100010_010;
      patterns[2012] = 19'b1010011000100010_010;
      patterns[2013] = 19'b1011011000100010_010;
      patterns[2014] = 19'b0100011000100000_110;
      patterns[2015] = 19'b1000011000100011_011;
      patterns[2016] = 19'b1001011000100011_011;
      patterns[2017] = 19'b1010011000100011_011;
      patterns[2018] = 19'b1011011000100011_011;
      patterns[2019] = 19'b0100011000100000_110;
      patterns[2020] = 19'b1000011000100100_100;
      patterns[2021] = 19'b1001011000100100_100;
      patterns[2022] = 19'b1010011000100100_100;
      patterns[2023] = 19'b1011011000100100_100;
      patterns[2024] = 19'b0100011000100000_110;
      patterns[2025] = 19'b1000011000100101_101;
      patterns[2026] = 19'b1001011000100101_101;
      patterns[2027] = 19'b1010011000100101_101;
      patterns[2028] = 19'b1011011000100101_101;
      patterns[2029] = 19'b0100011000100000_110;
      patterns[2030] = 19'b1000011000100110_110;
      patterns[2031] = 19'b1001011000100110_110;
      patterns[2032] = 19'b1010011000100110_110;
      patterns[2033] = 19'b1011011000100110_110;
      patterns[2034] = 19'b0100011000100000_110;
      patterns[2035] = 19'b1000011000100111_111;
      patterns[2036] = 19'b1001011000100111_111;
      patterns[2037] = 19'b1010011000100111_111;
      patterns[2038] = 19'b1011011000100111_111;
      patterns[2039] = 19'b0100011000100000_110;
      patterns[2040] = 19'b1000011000110000_000;
      patterns[2041] = 19'b1001011000110000_000;
      patterns[2042] = 19'b1010011000110000_000;
      patterns[2043] = 19'b1011011000110000_000;
      patterns[2044] = 19'b0100011000110000_110;
      patterns[2045] = 19'b1000011000110001_001;
      patterns[2046] = 19'b1001011000110001_001;
      patterns[2047] = 19'b1010011000110001_001;
      patterns[2048] = 19'b1011011000110001_001;
      patterns[2049] = 19'b0100011000110000_110;
      patterns[2050] = 19'b1000011000110010_010;
      patterns[2051] = 19'b1001011000110010_010;
      patterns[2052] = 19'b1010011000110010_010;
      patterns[2053] = 19'b1011011000110010_010;
      patterns[2054] = 19'b0100011000110000_110;
      patterns[2055] = 19'b1000011000110011_011;
      patterns[2056] = 19'b1001011000110011_011;
      patterns[2057] = 19'b1010011000110011_011;
      patterns[2058] = 19'b1011011000110011_011;
      patterns[2059] = 19'b0100011000110000_110;
      patterns[2060] = 19'b1000011000110100_100;
      patterns[2061] = 19'b1001011000110100_100;
      patterns[2062] = 19'b1010011000110100_100;
      patterns[2063] = 19'b1011011000110100_100;
      patterns[2064] = 19'b0100011000110000_110;
      patterns[2065] = 19'b1000011000110101_101;
      patterns[2066] = 19'b1001011000110101_101;
      patterns[2067] = 19'b1010011000110101_101;
      patterns[2068] = 19'b1011011000110101_101;
      patterns[2069] = 19'b0100011000110000_110;
      patterns[2070] = 19'b1000011000110110_110;
      patterns[2071] = 19'b1001011000110110_110;
      patterns[2072] = 19'b1010011000110110_110;
      patterns[2073] = 19'b1011011000110110_110;
      patterns[2074] = 19'b0100011000110000_110;
      patterns[2075] = 19'b1000011000110111_111;
      patterns[2076] = 19'b1001011000110111_111;
      patterns[2077] = 19'b1010011000110111_111;
      patterns[2078] = 19'b1011011000110111_111;
      patterns[2079] = 19'b0100011000110000_110;
      patterns[2080] = 19'b1000011001000000_000;
      patterns[2081] = 19'b1001011001000000_000;
      patterns[2082] = 19'b1010011001000000_000;
      patterns[2083] = 19'b1011011001000000_000;
      patterns[2084] = 19'b0100011001000000_110;
      patterns[2085] = 19'b1000011001000001_001;
      patterns[2086] = 19'b1001011001000001_001;
      patterns[2087] = 19'b1010011001000001_001;
      patterns[2088] = 19'b1011011001000001_001;
      patterns[2089] = 19'b0100011001000000_110;
      patterns[2090] = 19'b1000011001000010_010;
      patterns[2091] = 19'b1001011001000010_010;
      patterns[2092] = 19'b1010011001000010_010;
      patterns[2093] = 19'b1011011001000010_010;
      patterns[2094] = 19'b0100011001000000_110;
      patterns[2095] = 19'b1000011001000011_011;
      patterns[2096] = 19'b1001011001000011_011;
      patterns[2097] = 19'b1010011001000011_011;
      patterns[2098] = 19'b1011011001000011_011;
      patterns[2099] = 19'b0100011001000000_110;
      patterns[2100] = 19'b1000011001000100_100;
      patterns[2101] = 19'b1001011001000100_100;
      patterns[2102] = 19'b1010011001000100_100;
      patterns[2103] = 19'b1011011001000100_100;
      patterns[2104] = 19'b0100011001000000_110;
      patterns[2105] = 19'b1000011001000101_101;
      patterns[2106] = 19'b1001011001000101_101;
      patterns[2107] = 19'b1010011001000101_101;
      patterns[2108] = 19'b1011011001000101_101;
      patterns[2109] = 19'b0100011001000000_110;
      patterns[2110] = 19'b1000011001000110_110;
      patterns[2111] = 19'b1001011001000110_110;
      patterns[2112] = 19'b1010011001000110_110;
      patterns[2113] = 19'b1011011001000110_110;
      patterns[2114] = 19'b0100011001000000_110;
      patterns[2115] = 19'b1000011001000111_111;
      patterns[2116] = 19'b1001011001000111_111;
      patterns[2117] = 19'b1010011001000111_111;
      patterns[2118] = 19'b1011011001000111_111;
      patterns[2119] = 19'b0100011001000000_110;
      patterns[2120] = 19'b1000011001010000_000;
      patterns[2121] = 19'b1001011001010000_000;
      patterns[2122] = 19'b1010011001010000_000;
      patterns[2123] = 19'b1011011001010000_000;
      patterns[2124] = 19'b0100011001010000_110;
      patterns[2125] = 19'b1000011001010001_001;
      patterns[2126] = 19'b1001011001010001_001;
      patterns[2127] = 19'b1010011001010001_001;
      patterns[2128] = 19'b1011011001010001_001;
      patterns[2129] = 19'b0100011001010000_110;
      patterns[2130] = 19'b1000011001010010_010;
      patterns[2131] = 19'b1001011001010010_010;
      patterns[2132] = 19'b1010011001010010_010;
      patterns[2133] = 19'b1011011001010010_010;
      patterns[2134] = 19'b0100011001010000_110;
      patterns[2135] = 19'b1000011001010011_011;
      patterns[2136] = 19'b1001011001010011_011;
      patterns[2137] = 19'b1010011001010011_011;
      patterns[2138] = 19'b1011011001010011_011;
      patterns[2139] = 19'b0100011001010000_110;
      patterns[2140] = 19'b1000011001010100_100;
      patterns[2141] = 19'b1001011001010100_100;
      patterns[2142] = 19'b1010011001010100_100;
      patterns[2143] = 19'b1011011001010100_100;
      patterns[2144] = 19'b0100011001010000_110;
      patterns[2145] = 19'b1000011001010101_101;
      patterns[2146] = 19'b1001011001010101_101;
      patterns[2147] = 19'b1010011001010101_101;
      patterns[2148] = 19'b1011011001010101_101;
      patterns[2149] = 19'b0100011001010000_110;
      patterns[2150] = 19'b1000011001010110_110;
      patterns[2151] = 19'b1001011001010110_110;
      patterns[2152] = 19'b1010011001010110_110;
      patterns[2153] = 19'b1011011001010110_110;
      patterns[2154] = 19'b0100011001010000_110;
      patterns[2155] = 19'b1000011001010111_111;
      patterns[2156] = 19'b1001011001010111_111;
      patterns[2157] = 19'b1010011001010111_111;
      patterns[2158] = 19'b1011011001010111_111;
      patterns[2159] = 19'b0100011001010000_110;
      patterns[2160] = 19'b1000011001100000_000;
      patterns[2161] = 19'b1001011001100000_000;
      patterns[2162] = 19'b1010011001100000_000;
      patterns[2163] = 19'b1011011001100000_000;
      patterns[2164] = 19'b0100011001100000_110;
      patterns[2165] = 19'b1000011001100001_001;
      patterns[2166] = 19'b1001011001100001_001;
      patterns[2167] = 19'b1010011001100001_001;
      patterns[2168] = 19'b1011011001100001_001;
      patterns[2169] = 19'b0100011001100000_110;
      patterns[2170] = 19'b1000011001100010_010;
      patterns[2171] = 19'b1001011001100010_010;
      patterns[2172] = 19'b1010011001100010_010;
      patterns[2173] = 19'b1011011001100010_010;
      patterns[2174] = 19'b0100011001100000_110;
      patterns[2175] = 19'b1000011001100011_011;
      patterns[2176] = 19'b1001011001100011_011;
      patterns[2177] = 19'b1010011001100011_011;
      patterns[2178] = 19'b1011011001100011_011;
      patterns[2179] = 19'b0100011001100000_110;
      patterns[2180] = 19'b1000011001100100_100;
      patterns[2181] = 19'b1001011001100100_100;
      patterns[2182] = 19'b1010011001100100_100;
      patterns[2183] = 19'b1011011001100100_100;
      patterns[2184] = 19'b0100011001100000_110;
      patterns[2185] = 19'b1000011001100101_101;
      patterns[2186] = 19'b1001011001100101_101;
      patterns[2187] = 19'b1010011001100101_101;
      patterns[2188] = 19'b1011011001100101_101;
      patterns[2189] = 19'b0100011001100000_110;
      patterns[2190] = 19'b1000011001100110_110;
      patterns[2191] = 19'b1001011001100110_110;
      patterns[2192] = 19'b1010011001100110_110;
      patterns[2193] = 19'b1011011001100110_110;
      patterns[2194] = 19'b0100011001100000_110;
      patterns[2195] = 19'b1000011001100111_111;
      patterns[2196] = 19'b1001011001100111_111;
      patterns[2197] = 19'b1010011001100111_111;
      patterns[2198] = 19'b1011011001100111_111;
      patterns[2199] = 19'b0100011001100000_110;
      patterns[2200] = 19'b1000011001110000_000;
      patterns[2201] = 19'b1001011001110000_000;
      patterns[2202] = 19'b1010011001110000_000;
      patterns[2203] = 19'b1011011001110000_000;
      patterns[2204] = 19'b0100011001110000_110;
      patterns[2205] = 19'b1000011001110001_001;
      patterns[2206] = 19'b1001011001110001_001;
      patterns[2207] = 19'b1010011001110001_001;
      patterns[2208] = 19'b1011011001110001_001;
      patterns[2209] = 19'b0100011001110000_110;
      patterns[2210] = 19'b1000011001110010_010;
      patterns[2211] = 19'b1001011001110010_010;
      patterns[2212] = 19'b1010011001110010_010;
      patterns[2213] = 19'b1011011001110010_010;
      patterns[2214] = 19'b0100011001110000_110;
      patterns[2215] = 19'b1000011001110011_011;
      patterns[2216] = 19'b1001011001110011_011;
      patterns[2217] = 19'b1010011001110011_011;
      patterns[2218] = 19'b1011011001110011_011;
      patterns[2219] = 19'b0100011001110000_110;
      patterns[2220] = 19'b1000011001110100_100;
      patterns[2221] = 19'b1001011001110100_100;
      patterns[2222] = 19'b1010011001110100_100;
      patterns[2223] = 19'b1011011001110100_100;
      patterns[2224] = 19'b0100011001110000_110;
      patterns[2225] = 19'b1000011001110101_101;
      patterns[2226] = 19'b1001011001110101_101;
      patterns[2227] = 19'b1010011001110101_101;
      patterns[2228] = 19'b1011011001110101_101;
      patterns[2229] = 19'b0100011001110000_110;
      patterns[2230] = 19'b1000011001110110_110;
      patterns[2231] = 19'b1001011001110110_110;
      patterns[2232] = 19'b1010011001110110_110;
      patterns[2233] = 19'b1011011001110110_110;
      patterns[2234] = 19'b0100011001110000_110;
      patterns[2235] = 19'b1000011001110111_111;
      patterns[2236] = 19'b1001011001110111_111;
      patterns[2237] = 19'b1010011001110111_111;
      patterns[2238] = 19'b1011011001110111_111;
      patterns[2239] = 19'b0100011001110000_110;
      patterns[2240] = 19'b1000011100000000_000;
      patterns[2241] = 19'b1001011100000000_000;
      patterns[2242] = 19'b1010011100000000_000;
      patterns[2243] = 19'b1011011100000000_000;
      patterns[2244] = 19'b0100011100000000_111;
      patterns[2245] = 19'b1000011100000001_001;
      patterns[2246] = 19'b1001011100000001_001;
      patterns[2247] = 19'b1010011100000001_001;
      patterns[2248] = 19'b1011011100000001_001;
      patterns[2249] = 19'b0100011100000000_111;
      patterns[2250] = 19'b1000011100000010_010;
      patterns[2251] = 19'b1001011100000010_010;
      patterns[2252] = 19'b1010011100000010_010;
      patterns[2253] = 19'b1011011100000010_010;
      patterns[2254] = 19'b0100011100000000_111;
      patterns[2255] = 19'b1000011100000011_011;
      patterns[2256] = 19'b1001011100000011_011;
      patterns[2257] = 19'b1010011100000011_011;
      patterns[2258] = 19'b1011011100000011_011;
      patterns[2259] = 19'b0100011100000000_111;
      patterns[2260] = 19'b1000011100000100_100;
      patterns[2261] = 19'b1001011100000100_100;
      patterns[2262] = 19'b1010011100000100_100;
      patterns[2263] = 19'b1011011100000100_100;
      patterns[2264] = 19'b0100011100000000_111;
      patterns[2265] = 19'b1000011100000101_101;
      patterns[2266] = 19'b1001011100000101_101;
      patterns[2267] = 19'b1010011100000101_101;
      patterns[2268] = 19'b1011011100000101_101;
      patterns[2269] = 19'b0100011100000000_111;
      patterns[2270] = 19'b1000011100000110_110;
      patterns[2271] = 19'b1001011100000110_110;
      patterns[2272] = 19'b1010011100000110_110;
      patterns[2273] = 19'b1011011100000110_110;
      patterns[2274] = 19'b0100011100000000_111;
      patterns[2275] = 19'b1000011100000111_111;
      patterns[2276] = 19'b1001011100000111_111;
      patterns[2277] = 19'b1010011100000111_111;
      patterns[2278] = 19'b1011011100000111_111;
      patterns[2279] = 19'b0100011100000000_111;
      patterns[2280] = 19'b1000011100010000_000;
      patterns[2281] = 19'b1001011100010000_000;
      patterns[2282] = 19'b1010011100010000_000;
      patterns[2283] = 19'b1011011100010000_000;
      patterns[2284] = 19'b0100011100010000_111;
      patterns[2285] = 19'b1000011100010001_001;
      patterns[2286] = 19'b1001011100010001_001;
      patterns[2287] = 19'b1010011100010001_001;
      patterns[2288] = 19'b1011011100010001_001;
      patterns[2289] = 19'b0100011100010000_111;
      patterns[2290] = 19'b1000011100010010_010;
      patterns[2291] = 19'b1001011100010010_010;
      patterns[2292] = 19'b1010011100010010_010;
      patterns[2293] = 19'b1011011100010010_010;
      patterns[2294] = 19'b0100011100010000_111;
      patterns[2295] = 19'b1000011100010011_011;
      patterns[2296] = 19'b1001011100010011_011;
      patterns[2297] = 19'b1010011100010011_011;
      patterns[2298] = 19'b1011011100010011_011;
      patterns[2299] = 19'b0100011100010000_111;
      patterns[2300] = 19'b1000011100010100_100;
      patterns[2301] = 19'b1001011100010100_100;
      patterns[2302] = 19'b1010011100010100_100;
      patterns[2303] = 19'b1011011100010100_100;
      patterns[2304] = 19'b0100011100010000_111;
      patterns[2305] = 19'b1000011100010101_101;
      patterns[2306] = 19'b1001011100010101_101;
      patterns[2307] = 19'b1010011100010101_101;
      patterns[2308] = 19'b1011011100010101_101;
      patterns[2309] = 19'b0100011100010000_111;
      patterns[2310] = 19'b1000011100010110_110;
      patterns[2311] = 19'b1001011100010110_110;
      patterns[2312] = 19'b1010011100010110_110;
      patterns[2313] = 19'b1011011100010110_110;
      patterns[2314] = 19'b0100011100010000_111;
      patterns[2315] = 19'b1000011100010111_111;
      patterns[2316] = 19'b1001011100010111_111;
      patterns[2317] = 19'b1010011100010111_111;
      patterns[2318] = 19'b1011011100010111_111;
      patterns[2319] = 19'b0100011100010000_111;
      patterns[2320] = 19'b1000011100100000_000;
      patterns[2321] = 19'b1001011100100000_000;
      patterns[2322] = 19'b1010011100100000_000;
      patterns[2323] = 19'b1011011100100000_000;
      patterns[2324] = 19'b0100011100100000_111;
      patterns[2325] = 19'b1000011100100001_001;
      patterns[2326] = 19'b1001011100100001_001;
      patterns[2327] = 19'b1010011100100001_001;
      patterns[2328] = 19'b1011011100100001_001;
      patterns[2329] = 19'b0100011100100000_111;
      patterns[2330] = 19'b1000011100100010_010;
      patterns[2331] = 19'b1001011100100010_010;
      patterns[2332] = 19'b1010011100100010_010;
      patterns[2333] = 19'b1011011100100010_010;
      patterns[2334] = 19'b0100011100100000_111;
      patterns[2335] = 19'b1000011100100011_011;
      patterns[2336] = 19'b1001011100100011_011;
      patterns[2337] = 19'b1010011100100011_011;
      patterns[2338] = 19'b1011011100100011_011;
      patterns[2339] = 19'b0100011100100000_111;
      patterns[2340] = 19'b1000011100100100_100;
      patterns[2341] = 19'b1001011100100100_100;
      patterns[2342] = 19'b1010011100100100_100;
      patterns[2343] = 19'b1011011100100100_100;
      patterns[2344] = 19'b0100011100100000_111;
      patterns[2345] = 19'b1000011100100101_101;
      patterns[2346] = 19'b1001011100100101_101;
      patterns[2347] = 19'b1010011100100101_101;
      patterns[2348] = 19'b1011011100100101_101;
      patterns[2349] = 19'b0100011100100000_111;
      patterns[2350] = 19'b1000011100100110_110;
      patterns[2351] = 19'b1001011100100110_110;
      patterns[2352] = 19'b1010011100100110_110;
      patterns[2353] = 19'b1011011100100110_110;
      patterns[2354] = 19'b0100011100100000_111;
      patterns[2355] = 19'b1000011100100111_111;
      patterns[2356] = 19'b1001011100100111_111;
      patterns[2357] = 19'b1010011100100111_111;
      patterns[2358] = 19'b1011011100100111_111;
      patterns[2359] = 19'b0100011100100000_111;
      patterns[2360] = 19'b1000011100110000_000;
      patterns[2361] = 19'b1001011100110000_000;
      patterns[2362] = 19'b1010011100110000_000;
      patterns[2363] = 19'b1011011100110000_000;
      patterns[2364] = 19'b0100011100110000_111;
      patterns[2365] = 19'b1000011100110001_001;
      patterns[2366] = 19'b1001011100110001_001;
      patterns[2367] = 19'b1010011100110001_001;
      patterns[2368] = 19'b1011011100110001_001;
      patterns[2369] = 19'b0100011100110000_111;
      patterns[2370] = 19'b1000011100110010_010;
      patterns[2371] = 19'b1001011100110010_010;
      patterns[2372] = 19'b1010011100110010_010;
      patterns[2373] = 19'b1011011100110010_010;
      patterns[2374] = 19'b0100011100110000_111;
      patterns[2375] = 19'b1000011100110011_011;
      patterns[2376] = 19'b1001011100110011_011;
      patterns[2377] = 19'b1010011100110011_011;
      patterns[2378] = 19'b1011011100110011_011;
      patterns[2379] = 19'b0100011100110000_111;
      patterns[2380] = 19'b1000011100110100_100;
      patterns[2381] = 19'b1001011100110100_100;
      patterns[2382] = 19'b1010011100110100_100;
      patterns[2383] = 19'b1011011100110100_100;
      patterns[2384] = 19'b0100011100110000_111;
      patterns[2385] = 19'b1000011100110101_101;
      patterns[2386] = 19'b1001011100110101_101;
      patterns[2387] = 19'b1010011100110101_101;
      patterns[2388] = 19'b1011011100110101_101;
      patterns[2389] = 19'b0100011100110000_111;
      patterns[2390] = 19'b1000011100110110_110;
      patterns[2391] = 19'b1001011100110110_110;
      patterns[2392] = 19'b1010011100110110_110;
      patterns[2393] = 19'b1011011100110110_110;
      patterns[2394] = 19'b0100011100110000_111;
      patterns[2395] = 19'b1000011100110111_111;
      patterns[2396] = 19'b1001011100110111_111;
      patterns[2397] = 19'b1010011100110111_111;
      patterns[2398] = 19'b1011011100110111_111;
      patterns[2399] = 19'b0100011100110000_111;
      patterns[2400] = 19'b1000011101000000_000;
      patterns[2401] = 19'b1001011101000000_000;
      patterns[2402] = 19'b1010011101000000_000;
      patterns[2403] = 19'b1011011101000000_000;
      patterns[2404] = 19'b0100011101000000_111;
      patterns[2405] = 19'b1000011101000001_001;
      patterns[2406] = 19'b1001011101000001_001;
      patterns[2407] = 19'b1010011101000001_001;
      patterns[2408] = 19'b1011011101000001_001;
      patterns[2409] = 19'b0100011101000000_111;
      patterns[2410] = 19'b1000011101000010_010;
      patterns[2411] = 19'b1001011101000010_010;
      patterns[2412] = 19'b1010011101000010_010;
      patterns[2413] = 19'b1011011101000010_010;
      patterns[2414] = 19'b0100011101000000_111;
      patterns[2415] = 19'b1000011101000011_011;
      patterns[2416] = 19'b1001011101000011_011;
      patterns[2417] = 19'b1010011101000011_011;
      patterns[2418] = 19'b1011011101000011_011;
      patterns[2419] = 19'b0100011101000000_111;
      patterns[2420] = 19'b1000011101000100_100;
      patterns[2421] = 19'b1001011101000100_100;
      patterns[2422] = 19'b1010011101000100_100;
      patterns[2423] = 19'b1011011101000100_100;
      patterns[2424] = 19'b0100011101000000_111;
      patterns[2425] = 19'b1000011101000101_101;
      patterns[2426] = 19'b1001011101000101_101;
      patterns[2427] = 19'b1010011101000101_101;
      patterns[2428] = 19'b1011011101000101_101;
      patterns[2429] = 19'b0100011101000000_111;
      patterns[2430] = 19'b1000011101000110_110;
      patterns[2431] = 19'b1001011101000110_110;
      patterns[2432] = 19'b1010011101000110_110;
      patterns[2433] = 19'b1011011101000110_110;
      patterns[2434] = 19'b0100011101000000_111;
      patterns[2435] = 19'b1000011101000111_111;
      patterns[2436] = 19'b1001011101000111_111;
      patterns[2437] = 19'b1010011101000111_111;
      patterns[2438] = 19'b1011011101000111_111;
      patterns[2439] = 19'b0100011101000000_111;
      patterns[2440] = 19'b1000011101010000_000;
      patterns[2441] = 19'b1001011101010000_000;
      patterns[2442] = 19'b1010011101010000_000;
      patterns[2443] = 19'b1011011101010000_000;
      patterns[2444] = 19'b0100011101010000_111;
      patterns[2445] = 19'b1000011101010001_001;
      patterns[2446] = 19'b1001011101010001_001;
      patterns[2447] = 19'b1010011101010001_001;
      patterns[2448] = 19'b1011011101010001_001;
      patterns[2449] = 19'b0100011101010000_111;
      patterns[2450] = 19'b1000011101010010_010;
      patterns[2451] = 19'b1001011101010010_010;
      patterns[2452] = 19'b1010011101010010_010;
      patterns[2453] = 19'b1011011101010010_010;
      patterns[2454] = 19'b0100011101010000_111;
      patterns[2455] = 19'b1000011101010011_011;
      patterns[2456] = 19'b1001011101010011_011;
      patterns[2457] = 19'b1010011101010011_011;
      patterns[2458] = 19'b1011011101010011_011;
      patterns[2459] = 19'b0100011101010000_111;
      patterns[2460] = 19'b1000011101010100_100;
      patterns[2461] = 19'b1001011101010100_100;
      patterns[2462] = 19'b1010011101010100_100;
      patterns[2463] = 19'b1011011101010100_100;
      patterns[2464] = 19'b0100011101010000_111;
      patterns[2465] = 19'b1000011101010101_101;
      patterns[2466] = 19'b1001011101010101_101;
      patterns[2467] = 19'b1010011101010101_101;
      patterns[2468] = 19'b1011011101010101_101;
      patterns[2469] = 19'b0100011101010000_111;
      patterns[2470] = 19'b1000011101010110_110;
      patterns[2471] = 19'b1001011101010110_110;
      patterns[2472] = 19'b1010011101010110_110;
      patterns[2473] = 19'b1011011101010110_110;
      patterns[2474] = 19'b0100011101010000_111;
      patterns[2475] = 19'b1000011101010111_111;
      patterns[2476] = 19'b1001011101010111_111;
      patterns[2477] = 19'b1010011101010111_111;
      patterns[2478] = 19'b1011011101010111_111;
      patterns[2479] = 19'b0100011101010000_111;
      patterns[2480] = 19'b1000011101100000_000;
      patterns[2481] = 19'b1001011101100000_000;
      patterns[2482] = 19'b1010011101100000_000;
      patterns[2483] = 19'b1011011101100000_000;
      patterns[2484] = 19'b0100011101100000_111;
      patterns[2485] = 19'b1000011101100001_001;
      patterns[2486] = 19'b1001011101100001_001;
      patterns[2487] = 19'b1010011101100001_001;
      patterns[2488] = 19'b1011011101100001_001;
      patterns[2489] = 19'b0100011101100000_111;
      patterns[2490] = 19'b1000011101100010_010;
      patterns[2491] = 19'b1001011101100010_010;
      patterns[2492] = 19'b1010011101100010_010;
      patterns[2493] = 19'b1011011101100010_010;
      patterns[2494] = 19'b0100011101100000_111;
      patterns[2495] = 19'b1000011101100011_011;
      patterns[2496] = 19'b1001011101100011_011;
      patterns[2497] = 19'b1010011101100011_011;
      patterns[2498] = 19'b1011011101100011_011;
      patterns[2499] = 19'b0100011101100000_111;
      patterns[2500] = 19'b1000011101100100_100;
      patterns[2501] = 19'b1001011101100100_100;
      patterns[2502] = 19'b1010011101100100_100;
      patterns[2503] = 19'b1011011101100100_100;
      patterns[2504] = 19'b0100011101100000_111;
      patterns[2505] = 19'b1000011101100101_101;
      patterns[2506] = 19'b1001011101100101_101;
      patterns[2507] = 19'b1010011101100101_101;
      patterns[2508] = 19'b1011011101100101_101;
      patterns[2509] = 19'b0100011101100000_111;
      patterns[2510] = 19'b1000011101100110_110;
      patterns[2511] = 19'b1001011101100110_110;
      patterns[2512] = 19'b1010011101100110_110;
      patterns[2513] = 19'b1011011101100110_110;
      patterns[2514] = 19'b0100011101100000_111;
      patterns[2515] = 19'b1000011101100111_111;
      patterns[2516] = 19'b1001011101100111_111;
      patterns[2517] = 19'b1010011101100111_111;
      patterns[2518] = 19'b1011011101100111_111;
      patterns[2519] = 19'b0100011101100000_111;
      patterns[2520] = 19'b1000011101110000_000;
      patterns[2521] = 19'b1001011101110000_000;
      patterns[2522] = 19'b1010011101110000_000;
      patterns[2523] = 19'b1011011101110000_000;
      patterns[2524] = 19'b0100011101110000_111;
      patterns[2525] = 19'b1000011101110001_001;
      patterns[2526] = 19'b1001011101110001_001;
      patterns[2527] = 19'b1010011101110001_001;
      patterns[2528] = 19'b1011011101110001_001;
      patterns[2529] = 19'b0100011101110000_111;
      patterns[2530] = 19'b1000011101110010_010;
      patterns[2531] = 19'b1001011101110010_010;
      patterns[2532] = 19'b1010011101110010_010;
      patterns[2533] = 19'b1011011101110010_010;
      patterns[2534] = 19'b0100011101110000_111;
      patterns[2535] = 19'b1000011101110011_011;
      patterns[2536] = 19'b1001011101110011_011;
      patterns[2537] = 19'b1010011101110011_011;
      patterns[2538] = 19'b1011011101110011_011;
      patterns[2539] = 19'b0100011101110000_111;
      patterns[2540] = 19'b1000011101110100_100;
      patterns[2541] = 19'b1001011101110100_100;
      patterns[2542] = 19'b1010011101110100_100;
      patterns[2543] = 19'b1011011101110100_100;
      patterns[2544] = 19'b0100011101110000_111;
      patterns[2545] = 19'b1000011101110101_101;
      patterns[2546] = 19'b1001011101110101_101;
      patterns[2547] = 19'b1010011101110101_101;
      patterns[2548] = 19'b1011011101110101_101;
      patterns[2549] = 19'b0100011101110000_111;
      patterns[2550] = 19'b1000011101110110_110;
      patterns[2551] = 19'b1001011101110110_110;
      patterns[2552] = 19'b1010011101110110_110;
      patterns[2553] = 19'b1011011101110110_110;
      patterns[2554] = 19'b0100011101110000_111;
      patterns[2555] = 19'b1000011101110111_111;
      patterns[2556] = 19'b1001011101110111_111;
      patterns[2557] = 19'b1010011101110111_111;
      patterns[2558] = 19'b1011011101110111_111;
      patterns[2559] = 19'b0100011101110000_111;

      for (i = 0; i < 2560; i = i + 1)
      begin
        INST = patterns[i][18:3];
        #10;
        if (patterns[i][2:0] !== 3'hx)
        begin
          if (RS2 !== patterns[i][2:0])
          begin
            $display("%d:RS2: (assertion error). Expected %h, found %h", i, patterns[i][2:0], RS2);
            $finish;
          end
        end
      end

      $display("All tests passed.");
    end
    endmodule
