//  A testbench for control_unit_All Tests_tb
`timescale 1us/1ns

module control_unit_All Tests_tb;
    reg [15:0] INST;
    reg FL_Z;
    wire [1:0] ALUOP;
    wire [2:0] RS1;
    wire [2:0] RS2;
    wire [2:0] WS;
    wire STR;
    wire WE;
    wire [1:0] DMUX;
    wire LDR;
    wire FL_EN;
    wire HE;

  control_unit control_unit0 (
    .INST(INST),
    .FL_Z(FL_Z),
    .ALUOP(ALUOP),
    .RS1(RS1),
    .RS2(RS2),
    .WS(WS),
    .STR(STR),
    .WE(WE),
    .DMUX(DMUX),
    .LDR(LDR),
    .FL_EN(FL_EN),
    .HE(HE)
  );

    reg [32:0] patterns[0:10751];
    integer i;

    initial begin
      patterns[0] = 33'b1000000000000000_0_1_00_000_000_000_0_x_00;
      patterns[1] = 33'b1000100000000000_1_1_00_000_000_000_0_x_00;
      patterns[2] = 33'b1000100000000000_0_0_00_000_000_000_0_0_00;
      patterns[3] = 33'b1001000000000000_0_1_01_000_000_000_0_x_00;
      patterns[4] = 33'b1001100000000000_1_1_01_000_000_000_0_x_00;
      patterns[5] = 33'b1001100000000000_0_0_00_000_000_000_0_0_00;
      patterns[6] = 33'b1010000000000000_0_1_10_000_000_000_0_x_00;
      patterns[7] = 33'b1010100000000000_1_1_10_000_000_000_0_x_00;
      patterns[8] = 33'b1010100000000000_0_0_00_000_000_000_0_0_00;
      patterns[9] = 33'b1011000000000000_0_1_11_000_000_000_0_x_00;
      patterns[10] = 33'b1011100000000000_1_1_11_000_000_000_0_x_00;
      patterns[11] = 33'b1011100000000000_0_0_00_000_000_000_0_0_00;
      patterns[12] = 33'b0101000000000000_0_1_xx_000_xxx_000_0_1_01;
      patterns[13] = 33'b0101100000000000_1_1_xx_000_xxx_000_0_1_01;
      patterns[14] = 33'b0101100000000000_0_0_00_000_000_000_0_0_00;
      patterns[15] = 33'b0100000000000000_0_0_xx_000_000_xxx_1_x_xx;
      patterns[16] = 33'b0100100000000000_1_0_xx_000_000_xxx_1_x_xx;
      patterns[17] = 33'b0100100000000000_0_0_00_000_000_000_0_0_00;
      patterns[18] = 33'b0000000000001101_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[19] = 33'b0000100000001101_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[20] = 33'b0000100000001101_0_0_00_000_000_000_0_0_00;
      patterns[21] = 33'b1000000000000001_0_1_00_000_001_000_0_x_00;
      patterns[22] = 33'b1000100000000001_1_1_00_000_001_000_0_x_00;
      patterns[23] = 33'b1000100000000001_0_0_00_000_000_000_0_0_00;
      patterns[24] = 33'b1001000000000001_0_1_01_000_001_000_0_x_00;
      patterns[25] = 33'b1001100000000001_1_1_01_000_001_000_0_x_00;
      patterns[26] = 33'b1001100000000001_0_0_00_000_000_000_0_0_00;
      patterns[27] = 33'b1010000000000001_0_1_10_000_001_000_0_x_00;
      patterns[28] = 33'b1010100000000001_1_1_10_000_001_000_0_x_00;
      patterns[29] = 33'b1010100000000001_0_0_00_000_000_000_0_0_00;
      patterns[30] = 33'b1011000000000001_0_1_11_000_001_000_0_x_00;
      patterns[31] = 33'b1011100000000001_1_1_11_000_001_000_0_x_00;
      patterns[32] = 33'b1011100000000001_0_0_00_000_000_000_0_0_00;
      patterns[33] = 33'b0101000000000000_0_1_xx_000_xxx_000_0_1_01;
      patterns[34] = 33'b0101100000000000_1_1_xx_000_xxx_000_0_1_01;
      patterns[35] = 33'b0101100000000000_0_0_00_000_000_000_0_0_00;
      patterns[36] = 33'b0100000000000000_0_0_xx_000_000_xxx_1_x_xx;
      patterns[37] = 33'b0100100000000000_1_0_xx_000_000_xxx_1_x_xx;
      patterns[38] = 33'b0100100000000000_0_0_00_000_000_000_0_0_00;
      patterns[39] = 33'b0000000010010101_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[40] = 33'b0000100010010101_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[41] = 33'b0000100010010101_0_0_00_000_000_000_0_0_00;
      patterns[42] = 33'b1000000000000010_0_1_00_000_010_000_0_x_00;
      patterns[43] = 33'b1000100000000010_1_1_00_000_010_000_0_x_00;
      patterns[44] = 33'b1000100000000010_0_0_00_000_000_000_0_0_00;
      patterns[45] = 33'b1001000000000010_0_1_01_000_010_000_0_x_00;
      patterns[46] = 33'b1001100000000010_1_1_01_000_010_000_0_x_00;
      patterns[47] = 33'b1001100000000010_0_0_00_000_000_000_0_0_00;
      patterns[48] = 33'b1010000000000010_0_1_10_000_010_000_0_x_00;
      patterns[49] = 33'b1010100000000010_1_1_10_000_010_000_0_x_00;
      patterns[50] = 33'b1010100000000010_0_0_00_000_000_000_0_0_00;
      patterns[51] = 33'b1011000000000010_0_1_11_000_010_000_0_x_00;
      patterns[52] = 33'b1011100000000010_1_1_11_000_010_000_0_x_00;
      patterns[53] = 33'b1011100000000010_0_0_00_000_000_000_0_0_00;
      patterns[54] = 33'b0101000000000000_0_1_xx_000_xxx_000_0_1_01;
      patterns[55] = 33'b0101100000000000_1_1_xx_000_xxx_000_0_1_01;
      patterns[56] = 33'b0101100000000000_0_0_00_000_000_000_0_0_00;
      patterns[57] = 33'b0100000000000000_0_0_xx_000_000_xxx_1_x_xx;
      patterns[58] = 33'b0100100000000000_1_0_xx_000_000_xxx_1_x_xx;
      patterns[59] = 33'b0100100000000000_0_0_00_000_000_000_0_0_00;
      patterns[60] = 33'b0000000001000010_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[61] = 33'b0000100001000010_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[62] = 33'b0000100001000010_0_0_00_000_000_000_0_0_00;
      patterns[63] = 33'b1000000000000011_0_1_00_000_011_000_0_x_00;
      patterns[64] = 33'b1000100000000011_1_1_00_000_011_000_0_x_00;
      patterns[65] = 33'b1000100000000011_0_0_00_000_000_000_0_0_00;
      patterns[66] = 33'b1001000000000011_0_1_01_000_011_000_0_x_00;
      patterns[67] = 33'b1001100000000011_1_1_01_000_011_000_0_x_00;
      patterns[68] = 33'b1001100000000011_0_0_00_000_000_000_0_0_00;
      patterns[69] = 33'b1010000000000011_0_1_10_000_011_000_0_x_00;
      patterns[70] = 33'b1010100000000011_1_1_10_000_011_000_0_x_00;
      patterns[71] = 33'b1010100000000011_0_0_00_000_000_000_0_0_00;
      patterns[72] = 33'b1011000000000011_0_1_11_000_011_000_0_x_00;
      patterns[73] = 33'b1011100000000011_1_1_11_000_011_000_0_x_00;
      patterns[74] = 33'b1011100000000011_0_0_00_000_000_000_0_0_00;
      patterns[75] = 33'b0101000000000000_0_1_xx_000_xxx_000_0_1_01;
      patterns[76] = 33'b0101100000000000_1_1_xx_000_xxx_000_0_1_01;
      patterns[77] = 33'b0101100000000000_0_0_00_000_000_000_0_0_00;
      patterns[78] = 33'b0100000000000000_0_0_xx_000_000_xxx_1_x_xx;
      patterns[79] = 33'b0100100000000000_1_0_xx_000_000_xxx_1_x_xx;
      patterns[80] = 33'b0100100000000000_0_0_00_000_000_000_0_0_00;
      patterns[81] = 33'b0000000010110001_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[82] = 33'b0000100010110001_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[83] = 33'b0000100010110001_0_0_00_000_000_000_0_0_00;
      patterns[84] = 33'b1000000000000100_0_1_00_000_100_000_0_x_00;
      patterns[85] = 33'b1000100000000100_1_1_00_000_100_000_0_x_00;
      patterns[86] = 33'b1000100000000100_0_0_00_000_000_000_0_0_00;
      patterns[87] = 33'b1001000000000100_0_1_01_000_100_000_0_x_00;
      patterns[88] = 33'b1001100000000100_1_1_01_000_100_000_0_x_00;
      patterns[89] = 33'b1001100000000100_0_0_00_000_000_000_0_0_00;
      patterns[90] = 33'b1010000000000100_0_1_10_000_100_000_0_x_00;
      patterns[91] = 33'b1010100000000100_1_1_10_000_100_000_0_x_00;
      patterns[92] = 33'b1010100000000100_0_0_00_000_000_000_0_0_00;
      patterns[93] = 33'b1011000000000100_0_1_11_000_100_000_0_x_00;
      patterns[94] = 33'b1011100000000100_1_1_11_000_100_000_0_x_00;
      patterns[95] = 33'b1011100000000100_0_0_00_000_000_000_0_0_00;
      patterns[96] = 33'b0101000000000000_0_1_xx_000_xxx_000_0_1_01;
      patterns[97] = 33'b0101100000000000_1_1_xx_000_xxx_000_0_1_01;
      patterns[98] = 33'b0101100000000000_0_0_00_000_000_000_0_0_00;
      patterns[99] = 33'b0100000000000000_0_0_xx_000_000_xxx_1_x_xx;
      patterns[100] = 33'b0100100000000000_1_0_xx_000_000_xxx_1_x_xx;
      patterns[101] = 33'b0100100000000000_0_0_00_000_000_000_0_0_00;
      patterns[102] = 33'b0000000001110100_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[103] = 33'b0000100001110100_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[104] = 33'b0000100001110100_0_0_00_000_000_000_0_0_00;
      patterns[105] = 33'b1000000000000101_0_1_00_000_101_000_0_x_00;
      patterns[106] = 33'b1000100000000101_1_1_00_000_101_000_0_x_00;
      patterns[107] = 33'b1000100000000101_0_0_00_000_000_000_0_0_00;
      patterns[108] = 33'b1001000000000101_0_1_01_000_101_000_0_x_00;
      patterns[109] = 33'b1001100000000101_1_1_01_000_101_000_0_x_00;
      patterns[110] = 33'b1001100000000101_0_0_00_000_000_000_0_0_00;
      patterns[111] = 33'b1010000000000101_0_1_10_000_101_000_0_x_00;
      patterns[112] = 33'b1010100000000101_1_1_10_000_101_000_0_x_00;
      patterns[113] = 33'b1010100000000101_0_0_00_000_000_000_0_0_00;
      patterns[114] = 33'b1011000000000101_0_1_11_000_101_000_0_x_00;
      patterns[115] = 33'b1011100000000101_1_1_11_000_101_000_0_x_00;
      patterns[116] = 33'b1011100000000101_0_0_00_000_000_000_0_0_00;
      patterns[117] = 33'b0101000000000000_0_1_xx_000_xxx_000_0_1_01;
      patterns[118] = 33'b0101100000000000_1_1_xx_000_xxx_000_0_1_01;
      patterns[119] = 33'b0101100000000000_0_0_00_000_000_000_0_0_00;
      patterns[120] = 33'b0100000000000000_0_0_xx_000_000_xxx_1_x_xx;
      patterns[121] = 33'b0100100000000000_1_0_xx_000_000_xxx_1_x_xx;
      patterns[122] = 33'b0100100000000000_0_0_00_000_000_000_0_0_00;
      patterns[123] = 33'b0000000011001101_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[124] = 33'b0000100011001101_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[125] = 33'b0000100011001101_0_0_00_000_000_000_0_0_00;
      patterns[126] = 33'b1000000000000110_0_1_00_000_110_000_0_x_00;
      patterns[127] = 33'b1000100000000110_1_1_00_000_110_000_0_x_00;
      patterns[128] = 33'b1000100000000110_0_0_00_000_000_000_0_0_00;
      patterns[129] = 33'b1001000000000110_0_1_01_000_110_000_0_x_00;
      patterns[130] = 33'b1001100000000110_1_1_01_000_110_000_0_x_00;
      patterns[131] = 33'b1001100000000110_0_0_00_000_000_000_0_0_00;
      patterns[132] = 33'b1010000000000110_0_1_10_000_110_000_0_x_00;
      patterns[133] = 33'b1010100000000110_1_1_10_000_110_000_0_x_00;
      patterns[134] = 33'b1010100000000110_0_0_00_000_000_000_0_0_00;
      patterns[135] = 33'b1011000000000110_0_1_11_000_110_000_0_x_00;
      patterns[136] = 33'b1011100000000110_1_1_11_000_110_000_0_x_00;
      patterns[137] = 33'b1011100000000110_0_0_00_000_000_000_0_0_00;
      patterns[138] = 33'b0101000000000000_0_1_xx_000_xxx_000_0_1_01;
      patterns[139] = 33'b0101100000000000_1_1_xx_000_xxx_000_0_1_01;
      patterns[140] = 33'b0101100000000000_0_0_00_000_000_000_0_0_00;
      patterns[141] = 33'b0100000000000000_0_0_xx_000_000_xxx_1_x_xx;
      patterns[142] = 33'b0100100000000000_1_0_xx_000_000_xxx_1_x_xx;
      patterns[143] = 33'b0100100000000000_0_0_00_000_000_000_0_0_00;
      patterns[144] = 33'b0000000000110100_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[145] = 33'b0000100000110100_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[146] = 33'b0000100000110100_0_0_00_000_000_000_0_0_00;
      patterns[147] = 33'b1000000000000111_0_1_00_000_111_000_0_x_00;
      patterns[148] = 33'b1000100000000111_1_1_00_000_111_000_0_x_00;
      patterns[149] = 33'b1000100000000111_0_0_00_000_000_000_0_0_00;
      patterns[150] = 33'b1001000000000111_0_1_01_000_111_000_0_x_00;
      patterns[151] = 33'b1001100000000111_1_1_01_000_111_000_0_x_00;
      patterns[152] = 33'b1001100000000111_0_0_00_000_000_000_0_0_00;
      patterns[153] = 33'b1010000000000111_0_1_10_000_111_000_0_x_00;
      patterns[154] = 33'b1010100000000111_1_1_10_000_111_000_0_x_00;
      patterns[155] = 33'b1010100000000111_0_0_00_000_000_000_0_0_00;
      patterns[156] = 33'b1011000000000111_0_1_11_000_111_000_0_x_00;
      patterns[157] = 33'b1011100000000111_1_1_11_000_111_000_0_x_00;
      patterns[158] = 33'b1011100000000111_0_0_00_000_000_000_0_0_00;
      patterns[159] = 33'b0101000000000000_0_1_xx_000_xxx_000_0_1_01;
      patterns[160] = 33'b0101100000000000_1_1_xx_000_xxx_000_0_1_01;
      patterns[161] = 33'b0101100000000000_0_0_00_000_000_000_0_0_00;
      patterns[162] = 33'b0100000000000000_0_0_xx_000_000_xxx_1_x_xx;
      patterns[163] = 33'b0100100000000000_1_0_xx_000_000_xxx_1_x_xx;
      patterns[164] = 33'b0100100000000000_0_0_00_000_000_000_0_0_00;
      patterns[165] = 33'b0000000010110111_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[166] = 33'b0000100010110111_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[167] = 33'b0000100010110111_0_0_00_000_000_000_0_0_00;
      patterns[168] = 33'b1000000000010000_0_1_00_001_000_000_0_x_00;
      patterns[169] = 33'b1000100000010000_1_1_00_001_000_000_0_x_00;
      patterns[170] = 33'b1000100000010000_0_0_00_000_000_000_0_0_00;
      patterns[171] = 33'b1001000000010000_0_1_01_001_000_000_0_x_00;
      patterns[172] = 33'b1001100000010000_1_1_01_001_000_000_0_x_00;
      patterns[173] = 33'b1001100000010000_0_0_00_000_000_000_0_0_00;
      patterns[174] = 33'b1010000000010000_0_1_10_001_000_000_0_x_00;
      patterns[175] = 33'b1010100000010000_1_1_10_001_000_000_0_x_00;
      patterns[176] = 33'b1010100000010000_0_0_00_000_000_000_0_0_00;
      patterns[177] = 33'b1011000000010000_0_1_11_001_000_000_0_x_00;
      patterns[178] = 33'b1011100000010000_1_1_11_001_000_000_0_x_00;
      patterns[179] = 33'b1011100000010000_0_0_00_000_000_000_0_0_00;
      patterns[180] = 33'b0101000000010000_0_1_xx_001_xxx_000_0_1_01;
      patterns[181] = 33'b0101100000010000_1_1_xx_001_xxx_000_0_1_01;
      patterns[182] = 33'b0101100000010000_0_0_00_000_000_000_0_0_00;
      patterns[183] = 33'b0100000000010000_0_0_xx_001_000_xxx_1_x_xx;
      patterns[184] = 33'b0100100000010000_1_0_xx_001_000_xxx_1_x_xx;
      patterns[185] = 33'b0100100000010000_0_0_00_000_000_000_0_0_00;
      patterns[186] = 33'b0000000010011010_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[187] = 33'b0000100010011010_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[188] = 33'b0000100010011010_0_0_00_000_000_000_0_0_00;
      patterns[189] = 33'b1000000000010001_0_1_00_001_001_000_0_x_00;
      patterns[190] = 33'b1000100000010001_1_1_00_001_001_000_0_x_00;
      patterns[191] = 33'b1000100000010001_0_0_00_000_000_000_0_0_00;
      patterns[192] = 33'b1001000000010001_0_1_01_001_001_000_0_x_00;
      patterns[193] = 33'b1001100000010001_1_1_01_001_001_000_0_x_00;
      patterns[194] = 33'b1001100000010001_0_0_00_000_000_000_0_0_00;
      patterns[195] = 33'b1010000000010001_0_1_10_001_001_000_0_x_00;
      patterns[196] = 33'b1010100000010001_1_1_10_001_001_000_0_x_00;
      patterns[197] = 33'b1010100000010001_0_0_00_000_000_000_0_0_00;
      patterns[198] = 33'b1011000000010001_0_1_11_001_001_000_0_x_00;
      patterns[199] = 33'b1011100000010001_1_1_11_001_001_000_0_x_00;
      patterns[200] = 33'b1011100000010001_0_0_00_000_000_000_0_0_00;
      patterns[201] = 33'b0101000000010000_0_1_xx_001_xxx_000_0_1_01;
      patterns[202] = 33'b0101100000010000_1_1_xx_001_xxx_000_0_1_01;
      patterns[203] = 33'b0101100000010000_0_0_00_000_000_000_0_0_00;
      patterns[204] = 33'b0100000000010000_0_0_xx_001_000_xxx_1_x_xx;
      patterns[205] = 33'b0100100000010000_1_0_xx_001_000_xxx_1_x_xx;
      patterns[206] = 33'b0100100000010000_0_0_00_000_000_000_0_0_00;
      patterns[207] = 33'b0000000011110111_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[208] = 33'b0000100011110111_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[209] = 33'b0000100011110111_0_0_00_000_000_000_0_0_00;
      patterns[210] = 33'b1000000000010010_0_1_00_001_010_000_0_x_00;
      patterns[211] = 33'b1000100000010010_1_1_00_001_010_000_0_x_00;
      patterns[212] = 33'b1000100000010010_0_0_00_000_000_000_0_0_00;
      patterns[213] = 33'b1001000000010010_0_1_01_001_010_000_0_x_00;
      patterns[214] = 33'b1001100000010010_1_1_01_001_010_000_0_x_00;
      patterns[215] = 33'b1001100000010010_0_0_00_000_000_000_0_0_00;
      patterns[216] = 33'b1010000000010010_0_1_10_001_010_000_0_x_00;
      patterns[217] = 33'b1010100000010010_1_1_10_001_010_000_0_x_00;
      patterns[218] = 33'b1010100000010010_0_0_00_000_000_000_0_0_00;
      patterns[219] = 33'b1011000000010010_0_1_11_001_010_000_0_x_00;
      patterns[220] = 33'b1011100000010010_1_1_11_001_010_000_0_x_00;
      patterns[221] = 33'b1011100000010010_0_0_00_000_000_000_0_0_00;
      patterns[222] = 33'b0101000000010000_0_1_xx_001_xxx_000_0_1_01;
      patterns[223] = 33'b0101100000010000_1_1_xx_001_xxx_000_0_1_01;
      patterns[224] = 33'b0101100000010000_0_0_00_000_000_000_0_0_00;
      patterns[225] = 33'b0100000000010000_0_0_xx_001_000_xxx_1_x_xx;
      patterns[226] = 33'b0100100000010000_1_0_xx_001_000_xxx_1_x_xx;
      patterns[227] = 33'b0100100000010000_0_0_00_000_000_000_0_0_00;
      patterns[228] = 33'b0000000001001101_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[229] = 33'b0000100001001101_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[230] = 33'b0000100001001101_0_0_00_000_000_000_0_0_00;
      patterns[231] = 33'b1000000000010011_0_1_00_001_011_000_0_x_00;
      patterns[232] = 33'b1000100000010011_1_1_00_001_011_000_0_x_00;
      patterns[233] = 33'b1000100000010011_0_0_00_000_000_000_0_0_00;
      patterns[234] = 33'b1001000000010011_0_1_01_001_011_000_0_x_00;
      patterns[235] = 33'b1001100000010011_1_1_01_001_011_000_0_x_00;
      patterns[236] = 33'b1001100000010011_0_0_00_000_000_000_0_0_00;
      patterns[237] = 33'b1010000000010011_0_1_10_001_011_000_0_x_00;
      patterns[238] = 33'b1010100000010011_1_1_10_001_011_000_0_x_00;
      patterns[239] = 33'b1010100000010011_0_0_00_000_000_000_0_0_00;
      patterns[240] = 33'b1011000000010011_0_1_11_001_011_000_0_x_00;
      patterns[241] = 33'b1011100000010011_1_1_11_001_011_000_0_x_00;
      patterns[242] = 33'b1011100000010011_0_0_00_000_000_000_0_0_00;
      patterns[243] = 33'b0101000000010000_0_1_xx_001_xxx_000_0_1_01;
      patterns[244] = 33'b0101100000010000_1_1_xx_001_xxx_000_0_1_01;
      patterns[245] = 33'b0101100000010000_0_0_00_000_000_000_0_0_00;
      patterns[246] = 33'b0100000000010000_0_0_xx_001_000_xxx_1_x_xx;
      patterns[247] = 33'b0100100000010000_1_0_xx_001_000_xxx_1_x_xx;
      patterns[248] = 33'b0100100000010000_0_0_00_000_000_000_0_0_00;
      patterns[249] = 33'b0000000001000010_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[250] = 33'b0000100001000010_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[251] = 33'b0000100001000010_0_0_00_000_000_000_0_0_00;
      patterns[252] = 33'b1000000000010100_0_1_00_001_100_000_0_x_00;
      patterns[253] = 33'b1000100000010100_1_1_00_001_100_000_0_x_00;
      patterns[254] = 33'b1000100000010100_0_0_00_000_000_000_0_0_00;
      patterns[255] = 33'b1001000000010100_0_1_01_001_100_000_0_x_00;
      patterns[256] = 33'b1001100000010100_1_1_01_001_100_000_0_x_00;
      patterns[257] = 33'b1001100000010100_0_0_00_000_000_000_0_0_00;
      patterns[258] = 33'b1010000000010100_0_1_10_001_100_000_0_x_00;
      patterns[259] = 33'b1010100000010100_1_1_10_001_100_000_0_x_00;
      patterns[260] = 33'b1010100000010100_0_0_00_000_000_000_0_0_00;
      patterns[261] = 33'b1011000000010100_0_1_11_001_100_000_0_x_00;
      patterns[262] = 33'b1011100000010100_1_1_11_001_100_000_0_x_00;
      patterns[263] = 33'b1011100000010100_0_0_00_000_000_000_0_0_00;
      patterns[264] = 33'b0101000000010000_0_1_xx_001_xxx_000_0_1_01;
      patterns[265] = 33'b0101100000010000_1_1_xx_001_xxx_000_0_1_01;
      patterns[266] = 33'b0101100000010000_0_0_00_000_000_000_0_0_00;
      patterns[267] = 33'b0100000000010000_0_0_xx_001_000_xxx_1_x_xx;
      patterns[268] = 33'b0100100000010000_1_0_xx_001_000_xxx_1_x_xx;
      patterns[269] = 33'b0100100000010000_0_0_00_000_000_000_0_0_00;
      patterns[270] = 33'b0000000010010111_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[271] = 33'b0000100010010111_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[272] = 33'b0000100010010111_0_0_00_000_000_000_0_0_00;
      patterns[273] = 33'b1000000000010101_0_1_00_001_101_000_0_x_00;
      patterns[274] = 33'b1000100000010101_1_1_00_001_101_000_0_x_00;
      patterns[275] = 33'b1000100000010101_0_0_00_000_000_000_0_0_00;
      patterns[276] = 33'b1001000000010101_0_1_01_001_101_000_0_x_00;
      patterns[277] = 33'b1001100000010101_1_1_01_001_101_000_0_x_00;
      patterns[278] = 33'b1001100000010101_0_0_00_000_000_000_0_0_00;
      patterns[279] = 33'b1010000000010101_0_1_10_001_101_000_0_x_00;
      patterns[280] = 33'b1010100000010101_1_1_10_001_101_000_0_x_00;
      patterns[281] = 33'b1010100000010101_0_0_00_000_000_000_0_0_00;
      patterns[282] = 33'b1011000000010101_0_1_11_001_101_000_0_x_00;
      patterns[283] = 33'b1011100000010101_1_1_11_001_101_000_0_x_00;
      patterns[284] = 33'b1011100000010101_0_0_00_000_000_000_0_0_00;
      patterns[285] = 33'b0101000000010000_0_1_xx_001_xxx_000_0_1_01;
      patterns[286] = 33'b0101100000010000_1_1_xx_001_xxx_000_0_1_01;
      patterns[287] = 33'b0101100000010000_0_0_00_000_000_000_0_0_00;
      patterns[288] = 33'b0100000000010000_0_0_xx_001_000_xxx_1_x_xx;
      patterns[289] = 33'b0100100000010000_1_0_xx_001_000_xxx_1_x_xx;
      patterns[290] = 33'b0100100000010000_0_0_00_000_000_000_0_0_00;
      patterns[291] = 33'b0000000011001100_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[292] = 33'b0000100011001100_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[293] = 33'b0000100011001100_0_0_00_000_000_000_0_0_00;
      patterns[294] = 33'b1000000000010110_0_1_00_001_110_000_0_x_00;
      patterns[295] = 33'b1000100000010110_1_1_00_001_110_000_0_x_00;
      patterns[296] = 33'b1000100000010110_0_0_00_000_000_000_0_0_00;
      patterns[297] = 33'b1001000000010110_0_1_01_001_110_000_0_x_00;
      patterns[298] = 33'b1001100000010110_1_1_01_001_110_000_0_x_00;
      patterns[299] = 33'b1001100000010110_0_0_00_000_000_000_0_0_00;
      patterns[300] = 33'b1010000000010110_0_1_10_001_110_000_0_x_00;
      patterns[301] = 33'b1010100000010110_1_1_10_001_110_000_0_x_00;
      patterns[302] = 33'b1010100000010110_0_0_00_000_000_000_0_0_00;
      patterns[303] = 33'b1011000000010110_0_1_11_001_110_000_0_x_00;
      patterns[304] = 33'b1011100000010110_1_1_11_001_110_000_0_x_00;
      patterns[305] = 33'b1011100000010110_0_0_00_000_000_000_0_0_00;
      patterns[306] = 33'b0101000000010000_0_1_xx_001_xxx_000_0_1_01;
      patterns[307] = 33'b0101100000010000_1_1_xx_001_xxx_000_0_1_01;
      patterns[308] = 33'b0101100000010000_0_0_00_000_000_000_0_0_00;
      patterns[309] = 33'b0100000000010000_0_0_xx_001_000_xxx_1_x_xx;
      patterns[310] = 33'b0100100000010000_1_0_xx_001_000_xxx_1_x_xx;
      patterns[311] = 33'b0100100000010000_0_0_00_000_000_000_0_0_00;
      patterns[312] = 33'b0000000000100100_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[313] = 33'b0000100000100100_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[314] = 33'b0000100000100100_0_0_00_000_000_000_0_0_00;
      patterns[315] = 33'b1000000000010111_0_1_00_001_111_000_0_x_00;
      patterns[316] = 33'b1000100000010111_1_1_00_001_111_000_0_x_00;
      patterns[317] = 33'b1000100000010111_0_0_00_000_000_000_0_0_00;
      patterns[318] = 33'b1001000000010111_0_1_01_001_111_000_0_x_00;
      patterns[319] = 33'b1001100000010111_1_1_01_001_111_000_0_x_00;
      patterns[320] = 33'b1001100000010111_0_0_00_000_000_000_0_0_00;
      patterns[321] = 33'b1010000000010111_0_1_10_001_111_000_0_x_00;
      patterns[322] = 33'b1010100000010111_1_1_10_001_111_000_0_x_00;
      patterns[323] = 33'b1010100000010111_0_0_00_000_000_000_0_0_00;
      patterns[324] = 33'b1011000000010111_0_1_11_001_111_000_0_x_00;
      patterns[325] = 33'b1011100000010111_1_1_11_001_111_000_0_x_00;
      patterns[326] = 33'b1011100000010111_0_0_00_000_000_000_0_0_00;
      patterns[327] = 33'b0101000000010000_0_1_xx_001_xxx_000_0_1_01;
      patterns[328] = 33'b0101100000010000_1_1_xx_001_xxx_000_0_1_01;
      patterns[329] = 33'b0101100000010000_0_0_00_000_000_000_0_0_00;
      patterns[330] = 33'b0100000000010000_0_0_xx_001_000_xxx_1_x_xx;
      patterns[331] = 33'b0100100000010000_1_0_xx_001_000_xxx_1_x_xx;
      patterns[332] = 33'b0100100000010000_0_0_00_000_000_000_0_0_00;
      patterns[333] = 33'b0000000001100101_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[334] = 33'b0000100001100101_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[335] = 33'b0000100001100101_0_0_00_000_000_000_0_0_00;
      patterns[336] = 33'b1000000000100000_0_1_00_010_000_000_0_x_00;
      patterns[337] = 33'b1000100000100000_1_1_00_010_000_000_0_x_00;
      patterns[338] = 33'b1000100000100000_0_0_00_000_000_000_0_0_00;
      patterns[339] = 33'b1001000000100000_0_1_01_010_000_000_0_x_00;
      patterns[340] = 33'b1001100000100000_1_1_01_010_000_000_0_x_00;
      patterns[341] = 33'b1001100000100000_0_0_00_000_000_000_0_0_00;
      patterns[342] = 33'b1010000000100000_0_1_10_010_000_000_0_x_00;
      patterns[343] = 33'b1010100000100000_1_1_10_010_000_000_0_x_00;
      patterns[344] = 33'b1010100000100000_0_0_00_000_000_000_0_0_00;
      patterns[345] = 33'b1011000000100000_0_1_11_010_000_000_0_x_00;
      patterns[346] = 33'b1011100000100000_1_1_11_010_000_000_0_x_00;
      patterns[347] = 33'b1011100000100000_0_0_00_000_000_000_0_0_00;
      patterns[348] = 33'b0101000000100000_0_1_xx_010_xxx_000_0_1_01;
      patterns[349] = 33'b0101100000100000_1_1_xx_010_xxx_000_0_1_01;
      patterns[350] = 33'b0101100000100000_0_0_00_000_000_000_0_0_00;
      patterns[351] = 33'b0100000000100000_0_0_xx_010_000_xxx_1_x_xx;
      patterns[352] = 33'b0100100000100000_1_0_xx_010_000_xxx_1_x_xx;
      patterns[353] = 33'b0100100000100000_0_0_00_000_000_000_0_0_00;
      patterns[354] = 33'b0000000011110001_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[355] = 33'b0000100011110001_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[356] = 33'b0000100011110001_0_0_00_000_000_000_0_0_00;
      patterns[357] = 33'b1000000000100001_0_1_00_010_001_000_0_x_00;
      patterns[358] = 33'b1000100000100001_1_1_00_010_001_000_0_x_00;
      patterns[359] = 33'b1000100000100001_0_0_00_000_000_000_0_0_00;
      patterns[360] = 33'b1001000000100001_0_1_01_010_001_000_0_x_00;
      patterns[361] = 33'b1001100000100001_1_1_01_010_001_000_0_x_00;
      patterns[362] = 33'b1001100000100001_0_0_00_000_000_000_0_0_00;
      patterns[363] = 33'b1010000000100001_0_1_10_010_001_000_0_x_00;
      patterns[364] = 33'b1010100000100001_1_1_10_010_001_000_0_x_00;
      patterns[365] = 33'b1010100000100001_0_0_00_000_000_000_0_0_00;
      patterns[366] = 33'b1011000000100001_0_1_11_010_001_000_0_x_00;
      patterns[367] = 33'b1011100000100001_1_1_11_010_001_000_0_x_00;
      patterns[368] = 33'b1011100000100001_0_0_00_000_000_000_0_0_00;
      patterns[369] = 33'b0101000000100000_0_1_xx_010_xxx_000_0_1_01;
      patterns[370] = 33'b0101100000100000_1_1_xx_010_xxx_000_0_1_01;
      patterns[371] = 33'b0101100000100000_0_0_00_000_000_000_0_0_00;
      patterns[372] = 33'b0100000000100000_0_0_xx_010_000_xxx_1_x_xx;
      patterns[373] = 33'b0100100000100000_1_0_xx_010_000_xxx_1_x_xx;
      patterns[374] = 33'b0100100000100000_0_0_00_000_000_000_0_0_00;
      patterns[375] = 33'b0000000001010110_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[376] = 33'b0000100001010110_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[377] = 33'b0000100001010110_0_0_00_000_000_000_0_0_00;
      patterns[378] = 33'b1000000000100010_0_1_00_010_010_000_0_x_00;
      patterns[379] = 33'b1000100000100010_1_1_00_010_010_000_0_x_00;
      patterns[380] = 33'b1000100000100010_0_0_00_000_000_000_0_0_00;
      patterns[381] = 33'b1001000000100010_0_1_01_010_010_000_0_x_00;
      patterns[382] = 33'b1001100000100010_1_1_01_010_010_000_0_x_00;
      patterns[383] = 33'b1001100000100010_0_0_00_000_000_000_0_0_00;
      patterns[384] = 33'b1010000000100010_0_1_10_010_010_000_0_x_00;
      patterns[385] = 33'b1010100000100010_1_1_10_010_010_000_0_x_00;
      patterns[386] = 33'b1010100000100010_0_0_00_000_000_000_0_0_00;
      patterns[387] = 33'b1011000000100010_0_1_11_010_010_000_0_x_00;
      patterns[388] = 33'b1011100000100010_1_1_11_010_010_000_0_x_00;
      patterns[389] = 33'b1011100000100010_0_0_00_000_000_000_0_0_00;
      patterns[390] = 33'b0101000000100000_0_1_xx_010_xxx_000_0_1_01;
      patterns[391] = 33'b0101100000100000_1_1_xx_010_xxx_000_0_1_01;
      patterns[392] = 33'b0101100000100000_0_0_00_000_000_000_0_0_00;
      patterns[393] = 33'b0100000000100000_0_0_xx_010_000_xxx_1_x_xx;
      patterns[394] = 33'b0100100000100000_1_0_xx_010_000_xxx_1_x_xx;
      patterns[395] = 33'b0100100000100000_0_0_00_000_000_000_0_0_00;
      patterns[396] = 33'b0000000000101000_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[397] = 33'b0000100000101000_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[398] = 33'b0000100000101000_0_0_00_000_000_000_0_0_00;
      patterns[399] = 33'b1000000000100011_0_1_00_010_011_000_0_x_00;
      patterns[400] = 33'b1000100000100011_1_1_00_010_011_000_0_x_00;
      patterns[401] = 33'b1000100000100011_0_0_00_000_000_000_0_0_00;
      patterns[402] = 33'b1001000000100011_0_1_01_010_011_000_0_x_00;
      patterns[403] = 33'b1001100000100011_1_1_01_010_011_000_0_x_00;
      patterns[404] = 33'b1001100000100011_0_0_00_000_000_000_0_0_00;
      patterns[405] = 33'b1010000000100011_0_1_10_010_011_000_0_x_00;
      patterns[406] = 33'b1010100000100011_1_1_10_010_011_000_0_x_00;
      patterns[407] = 33'b1010100000100011_0_0_00_000_000_000_0_0_00;
      patterns[408] = 33'b1011000000100011_0_1_11_010_011_000_0_x_00;
      patterns[409] = 33'b1011100000100011_1_1_11_010_011_000_0_x_00;
      patterns[410] = 33'b1011100000100011_0_0_00_000_000_000_0_0_00;
      patterns[411] = 33'b0101000000100000_0_1_xx_010_xxx_000_0_1_01;
      patterns[412] = 33'b0101100000100000_1_1_xx_010_xxx_000_0_1_01;
      patterns[413] = 33'b0101100000100000_0_0_00_000_000_000_0_0_00;
      patterns[414] = 33'b0100000000100000_0_0_xx_010_000_xxx_1_x_xx;
      patterns[415] = 33'b0100100000100000_1_0_xx_010_000_xxx_1_x_xx;
      patterns[416] = 33'b0100100000100000_0_0_00_000_000_000_0_0_00;
      patterns[417] = 33'b0000000001001001_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[418] = 33'b0000100001001001_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[419] = 33'b0000100001001001_0_0_00_000_000_000_0_0_00;
      patterns[420] = 33'b1000000000100100_0_1_00_010_100_000_0_x_00;
      patterns[421] = 33'b1000100000100100_1_1_00_010_100_000_0_x_00;
      patterns[422] = 33'b1000100000100100_0_0_00_000_000_000_0_0_00;
      patterns[423] = 33'b1001000000100100_0_1_01_010_100_000_0_x_00;
      patterns[424] = 33'b1001100000100100_1_1_01_010_100_000_0_x_00;
      patterns[425] = 33'b1001100000100100_0_0_00_000_000_000_0_0_00;
      patterns[426] = 33'b1010000000100100_0_1_10_010_100_000_0_x_00;
      patterns[427] = 33'b1010100000100100_1_1_10_010_100_000_0_x_00;
      patterns[428] = 33'b1010100000100100_0_0_00_000_000_000_0_0_00;
      patterns[429] = 33'b1011000000100100_0_1_11_010_100_000_0_x_00;
      patterns[430] = 33'b1011100000100100_1_1_11_010_100_000_0_x_00;
      patterns[431] = 33'b1011100000100100_0_0_00_000_000_000_0_0_00;
      patterns[432] = 33'b0101000000100000_0_1_xx_010_xxx_000_0_1_01;
      patterns[433] = 33'b0101100000100000_1_1_xx_010_xxx_000_0_1_01;
      patterns[434] = 33'b0101100000100000_0_0_00_000_000_000_0_0_00;
      patterns[435] = 33'b0100000000100000_0_0_xx_010_000_xxx_1_x_xx;
      patterns[436] = 33'b0100100000100000_1_0_xx_010_000_xxx_1_x_xx;
      patterns[437] = 33'b0100100000100000_0_0_00_000_000_000_0_0_00;
      patterns[438] = 33'b0000000001000011_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[439] = 33'b0000100001000011_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[440] = 33'b0000100001000011_0_0_00_000_000_000_0_0_00;
      patterns[441] = 33'b1000000000100101_0_1_00_010_101_000_0_x_00;
      patterns[442] = 33'b1000100000100101_1_1_00_010_101_000_0_x_00;
      patterns[443] = 33'b1000100000100101_0_0_00_000_000_000_0_0_00;
      patterns[444] = 33'b1001000000100101_0_1_01_010_101_000_0_x_00;
      patterns[445] = 33'b1001100000100101_1_1_01_010_101_000_0_x_00;
      patterns[446] = 33'b1001100000100101_0_0_00_000_000_000_0_0_00;
      patterns[447] = 33'b1010000000100101_0_1_10_010_101_000_0_x_00;
      patterns[448] = 33'b1010100000100101_1_1_10_010_101_000_0_x_00;
      patterns[449] = 33'b1010100000100101_0_0_00_000_000_000_0_0_00;
      patterns[450] = 33'b1011000000100101_0_1_11_010_101_000_0_x_00;
      patterns[451] = 33'b1011100000100101_1_1_11_010_101_000_0_x_00;
      patterns[452] = 33'b1011100000100101_0_0_00_000_000_000_0_0_00;
      patterns[453] = 33'b0101000000100000_0_1_xx_010_xxx_000_0_1_01;
      patterns[454] = 33'b0101100000100000_1_1_xx_010_xxx_000_0_1_01;
      patterns[455] = 33'b0101100000100000_0_0_00_000_000_000_0_0_00;
      patterns[456] = 33'b0100000000100000_0_0_xx_010_000_xxx_1_x_xx;
      patterns[457] = 33'b0100100000100000_1_0_xx_010_000_xxx_1_x_xx;
      patterns[458] = 33'b0100100000100000_0_0_00_000_000_000_0_0_00;
      patterns[459] = 33'b0000000010010011_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[460] = 33'b0000100010010011_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[461] = 33'b0000100010010011_0_0_00_000_000_000_0_0_00;
      patterns[462] = 33'b1000000000100110_0_1_00_010_110_000_0_x_00;
      patterns[463] = 33'b1000100000100110_1_1_00_010_110_000_0_x_00;
      patterns[464] = 33'b1000100000100110_0_0_00_000_000_000_0_0_00;
      patterns[465] = 33'b1001000000100110_0_1_01_010_110_000_0_x_00;
      patterns[466] = 33'b1001100000100110_1_1_01_010_110_000_0_x_00;
      patterns[467] = 33'b1001100000100110_0_0_00_000_000_000_0_0_00;
      patterns[468] = 33'b1010000000100110_0_1_10_010_110_000_0_x_00;
      patterns[469] = 33'b1010100000100110_1_1_10_010_110_000_0_x_00;
      patterns[470] = 33'b1010100000100110_0_0_00_000_000_000_0_0_00;
      patterns[471] = 33'b1011000000100110_0_1_11_010_110_000_0_x_00;
      patterns[472] = 33'b1011100000100110_1_1_11_010_110_000_0_x_00;
      patterns[473] = 33'b1011100000100110_0_0_00_000_000_000_0_0_00;
      patterns[474] = 33'b0101000000100000_0_1_xx_010_xxx_000_0_1_01;
      patterns[475] = 33'b0101100000100000_1_1_xx_010_xxx_000_0_1_01;
      patterns[476] = 33'b0101100000100000_0_0_00_000_000_000_0_0_00;
      patterns[477] = 33'b0100000000100000_0_0_xx_010_000_xxx_1_x_xx;
      patterns[478] = 33'b0100100000100000_1_0_xx_010_000_xxx_1_x_xx;
      patterns[479] = 33'b0100100000100000_0_0_00_000_000_000_0_0_00;
      patterns[480] = 33'b0000000010010111_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[481] = 33'b0000100010010111_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[482] = 33'b0000100010010111_0_0_00_000_000_000_0_0_00;
      patterns[483] = 33'b1000000000100111_0_1_00_010_111_000_0_x_00;
      patterns[484] = 33'b1000100000100111_1_1_00_010_111_000_0_x_00;
      patterns[485] = 33'b1000100000100111_0_0_00_000_000_000_0_0_00;
      patterns[486] = 33'b1001000000100111_0_1_01_010_111_000_0_x_00;
      patterns[487] = 33'b1001100000100111_1_1_01_010_111_000_0_x_00;
      patterns[488] = 33'b1001100000100111_0_0_00_000_000_000_0_0_00;
      patterns[489] = 33'b1010000000100111_0_1_10_010_111_000_0_x_00;
      patterns[490] = 33'b1010100000100111_1_1_10_010_111_000_0_x_00;
      patterns[491] = 33'b1010100000100111_0_0_00_000_000_000_0_0_00;
      patterns[492] = 33'b1011000000100111_0_1_11_010_111_000_0_x_00;
      patterns[493] = 33'b1011100000100111_1_1_11_010_111_000_0_x_00;
      patterns[494] = 33'b1011100000100111_0_0_00_000_000_000_0_0_00;
      patterns[495] = 33'b0101000000100000_0_1_xx_010_xxx_000_0_1_01;
      patterns[496] = 33'b0101100000100000_1_1_xx_010_xxx_000_0_1_01;
      patterns[497] = 33'b0101100000100000_0_0_00_000_000_000_0_0_00;
      patterns[498] = 33'b0100000000100000_0_0_xx_010_000_xxx_1_x_xx;
      patterns[499] = 33'b0100100000100000_1_0_xx_010_000_xxx_1_x_xx;
      patterns[500] = 33'b0100100000100000_0_0_00_000_000_000_0_0_00;
      patterns[501] = 33'b0000000000100100_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[502] = 33'b0000100000100100_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[503] = 33'b0000100000100100_0_0_00_000_000_000_0_0_00;
      patterns[504] = 33'b1000000000110000_0_1_00_011_000_000_0_x_00;
      patterns[505] = 33'b1000100000110000_1_1_00_011_000_000_0_x_00;
      patterns[506] = 33'b1000100000110000_0_0_00_000_000_000_0_0_00;
      patterns[507] = 33'b1001000000110000_0_1_01_011_000_000_0_x_00;
      patterns[508] = 33'b1001100000110000_1_1_01_011_000_000_0_x_00;
      patterns[509] = 33'b1001100000110000_0_0_00_000_000_000_0_0_00;
      patterns[510] = 33'b1010000000110000_0_1_10_011_000_000_0_x_00;
      patterns[511] = 33'b1010100000110000_1_1_10_011_000_000_0_x_00;
      patterns[512] = 33'b1010100000110000_0_0_00_000_000_000_0_0_00;
      patterns[513] = 33'b1011000000110000_0_1_11_011_000_000_0_x_00;
      patterns[514] = 33'b1011100000110000_1_1_11_011_000_000_0_x_00;
      patterns[515] = 33'b1011100000110000_0_0_00_000_000_000_0_0_00;
      patterns[516] = 33'b0101000000110000_0_1_xx_011_xxx_000_0_1_01;
      patterns[517] = 33'b0101100000110000_1_1_xx_011_xxx_000_0_1_01;
      patterns[518] = 33'b0101100000110000_0_0_00_000_000_000_0_0_00;
      patterns[519] = 33'b0100000000110000_0_0_xx_011_000_xxx_1_x_xx;
      patterns[520] = 33'b0100100000110000_1_0_xx_011_000_xxx_1_x_xx;
      patterns[521] = 33'b0100100000110000_0_0_00_000_000_000_0_0_00;
      patterns[522] = 33'b0000000001001000_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[523] = 33'b0000100001001000_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[524] = 33'b0000100001001000_0_0_00_000_000_000_0_0_00;
      patterns[525] = 33'b1000000000110001_0_1_00_011_001_000_0_x_00;
      patterns[526] = 33'b1000100000110001_1_1_00_011_001_000_0_x_00;
      patterns[527] = 33'b1000100000110001_0_0_00_000_000_000_0_0_00;
      patterns[528] = 33'b1001000000110001_0_1_01_011_001_000_0_x_00;
      patterns[529] = 33'b1001100000110001_1_1_01_011_001_000_0_x_00;
      patterns[530] = 33'b1001100000110001_0_0_00_000_000_000_0_0_00;
      patterns[531] = 33'b1010000000110001_0_1_10_011_001_000_0_x_00;
      patterns[532] = 33'b1010100000110001_1_1_10_011_001_000_0_x_00;
      patterns[533] = 33'b1010100000110001_0_0_00_000_000_000_0_0_00;
      patterns[534] = 33'b1011000000110001_0_1_11_011_001_000_0_x_00;
      patterns[535] = 33'b1011100000110001_1_1_11_011_001_000_0_x_00;
      patterns[536] = 33'b1011100000110001_0_0_00_000_000_000_0_0_00;
      patterns[537] = 33'b0101000000110000_0_1_xx_011_xxx_000_0_1_01;
      patterns[538] = 33'b0101100000110000_1_1_xx_011_xxx_000_0_1_01;
      patterns[539] = 33'b0101100000110000_0_0_00_000_000_000_0_0_00;
      patterns[540] = 33'b0100000000110000_0_0_xx_011_000_xxx_1_x_xx;
      patterns[541] = 33'b0100100000110000_1_0_xx_011_000_xxx_1_x_xx;
      patterns[542] = 33'b0100100000110000_0_0_00_000_000_000_0_0_00;
      patterns[543] = 33'b0000000010100110_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[544] = 33'b0000100010100110_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[545] = 33'b0000100010100110_0_0_00_000_000_000_0_0_00;
      patterns[546] = 33'b1000000000110010_0_1_00_011_010_000_0_x_00;
      patterns[547] = 33'b1000100000110010_1_1_00_011_010_000_0_x_00;
      patterns[548] = 33'b1000100000110010_0_0_00_000_000_000_0_0_00;
      patterns[549] = 33'b1001000000110010_0_1_01_011_010_000_0_x_00;
      patterns[550] = 33'b1001100000110010_1_1_01_011_010_000_0_x_00;
      patterns[551] = 33'b1001100000110010_0_0_00_000_000_000_0_0_00;
      patterns[552] = 33'b1010000000110010_0_1_10_011_010_000_0_x_00;
      patterns[553] = 33'b1010100000110010_1_1_10_011_010_000_0_x_00;
      patterns[554] = 33'b1010100000110010_0_0_00_000_000_000_0_0_00;
      patterns[555] = 33'b1011000000110010_0_1_11_011_010_000_0_x_00;
      patterns[556] = 33'b1011100000110010_1_1_11_011_010_000_0_x_00;
      patterns[557] = 33'b1011100000110010_0_0_00_000_000_000_0_0_00;
      patterns[558] = 33'b0101000000110000_0_1_xx_011_xxx_000_0_1_01;
      patterns[559] = 33'b0101100000110000_1_1_xx_011_xxx_000_0_1_01;
      patterns[560] = 33'b0101100000110000_0_0_00_000_000_000_0_0_00;
      patterns[561] = 33'b0100000000110000_0_0_xx_011_000_xxx_1_x_xx;
      patterns[562] = 33'b0100100000110000_1_0_xx_011_000_xxx_1_x_xx;
      patterns[563] = 33'b0100100000110000_0_0_00_000_000_000_0_0_00;
      patterns[564] = 33'b0000000010111101_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[565] = 33'b0000100010111101_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[566] = 33'b0000100010111101_0_0_00_000_000_000_0_0_00;
      patterns[567] = 33'b1000000000110011_0_1_00_011_011_000_0_x_00;
      patterns[568] = 33'b1000100000110011_1_1_00_011_011_000_0_x_00;
      patterns[569] = 33'b1000100000110011_0_0_00_000_000_000_0_0_00;
      patterns[570] = 33'b1001000000110011_0_1_01_011_011_000_0_x_00;
      patterns[571] = 33'b1001100000110011_1_1_01_011_011_000_0_x_00;
      patterns[572] = 33'b1001100000110011_0_0_00_000_000_000_0_0_00;
      patterns[573] = 33'b1010000000110011_0_1_10_011_011_000_0_x_00;
      patterns[574] = 33'b1010100000110011_1_1_10_011_011_000_0_x_00;
      patterns[575] = 33'b1010100000110011_0_0_00_000_000_000_0_0_00;
      patterns[576] = 33'b1011000000110011_0_1_11_011_011_000_0_x_00;
      patterns[577] = 33'b1011100000110011_1_1_11_011_011_000_0_x_00;
      patterns[578] = 33'b1011100000110011_0_0_00_000_000_000_0_0_00;
      patterns[579] = 33'b0101000000110000_0_1_xx_011_xxx_000_0_1_01;
      patterns[580] = 33'b0101100000110000_1_1_xx_011_xxx_000_0_1_01;
      patterns[581] = 33'b0101100000110000_0_0_00_000_000_000_0_0_00;
      patterns[582] = 33'b0100000000110000_0_0_xx_011_000_xxx_1_x_xx;
      patterns[583] = 33'b0100100000110000_1_0_xx_011_000_xxx_1_x_xx;
      patterns[584] = 33'b0100100000110000_0_0_00_000_000_000_0_0_00;
      patterns[585] = 33'b0000000001011110_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[586] = 33'b0000100001011110_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[587] = 33'b0000100001011110_0_0_00_000_000_000_0_0_00;
      patterns[588] = 33'b1000000000110100_0_1_00_011_100_000_0_x_00;
      patterns[589] = 33'b1000100000110100_1_1_00_011_100_000_0_x_00;
      patterns[590] = 33'b1000100000110100_0_0_00_000_000_000_0_0_00;
      patterns[591] = 33'b1001000000110100_0_1_01_011_100_000_0_x_00;
      patterns[592] = 33'b1001100000110100_1_1_01_011_100_000_0_x_00;
      patterns[593] = 33'b1001100000110100_0_0_00_000_000_000_0_0_00;
      patterns[594] = 33'b1010000000110100_0_1_10_011_100_000_0_x_00;
      patterns[595] = 33'b1010100000110100_1_1_10_011_100_000_0_x_00;
      patterns[596] = 33'b1010100000110100_0_0_00_000_000_000_0_0_00;
      patterns[597] = 33'b1011000000110100_0_1_11_011_100_000_0_x_00;
      patterns[598] = 33'b1011100000110100_1_1_11_011_100_000_0_x_00;
      patterns[599] = 33'b1011100000110100_0_0_00_000_000_000_0_0_00;
      patterns[600] = 33'b0101000000110000_0_1_xx_011_xxx_000_0_1_01;
      patterns[601] = 33'b0101100000110000_1_1_xx_011_xxx_000_0_1_01;
      patterns[602] = 33'b0101100000110000_0_0_00_000_000_000_0_0_00;
      patterns[603] = 33'b0100000000110000_0_0_xx_011_000_xxx_1_x_xx;
      patterns[604] = 33'b0100100000110000_1_0_xx_011_000_xxx_1_x_xx;
      patterns[605] = 33'b0100100000110000_0_0_00_000_000_000_0_0_00;
      patterns[606] = 33'b0000000011110110_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[607] = 33'b0000100011110110_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[608] = 33'b0000100011110110_0_0_00_000_000_000_0_0_00;
      patterns[609] = 33'b1000000000110101_0_1_00_011_101_000_0_x_00;
      patterns[610] = 33'b1000100000110101_1_1_00_011_101_000_0_x_00;
      patterns[611] = 33'b1000100000110101_0_0_00_000_000_000_0_0_00;
      patterns[612] = 33'b1001000000110101_0_1_01_011_101_000_0_x_00;
      patterns[613] = 33'b1001100000110101_1_1_01_011_101_000_0_x_00;
      patterns[614] = 33'b1001100000110101_0_0_00_000_000_000_0_0_00;
      patterns[615] = 33'b1010000000110101_0_1_10_011_101_000_0_x_00;
      patterns[616] = 33'b1010100000110101_1_1_10_011_101_000_0_x_00;
      patterns[617] = 33'b1010100000110101_0_0_00_000_000_000_0_0_00;
      patterns[618] = 33'b1011000000110101_0_1_11_011_101_000_0_x_00;
      patterns[619] = 33'b1011100000110101_1_1_11_011_101_000_0_x_00;
      patterns[620] = 33'b1011100000110101_0_0_00_000_000_000_0_0_00;
      patterns[621] = 33'b0101000000110000_0_1_xx_011_xxx_000_0_1_01;
      patterns[622] = 33'b0101100000110000_1_1_xx_011_xxx_000_0_1_01;
      patterns[623] = 33'b0101100000110000_0_0_00_000_000_000_0_0_00;
      patterns[624] = 33'b0100000000110000_0_0_xx_011_000_xxx_1_x_xx;
      patterns[625] = 33'b0100100000110000_1_0_xx_011_000_xxx_1_x_xx;
      patterns[626] = 33'b0100100000110000_0_0_00_000_000_000_0_0_00;
      patterns[627] = 33'b0000000001000000_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[628] = 33'b0000100001000000_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[629] = 33'b0000100001000000_0_0_00_000_000_000_0_0_00;
      patterns[630] = 33'b1000000000110110_0_1_00_011_110_000_0_x_00;
      patterns[631] = 33'b1000100000110110_1_1_00_011_110_000_0_x_00;
      patterns[632] = 33'b1000100000110110_0_0_00_000_000_000_0_0_00;
      patterns[633] = 33'b1001000000110110_0_1_01_011_110_000_0_x_00;
      patterns[634] = 33'b1001100000110110_1_1_01_011_110_000_0_x_00;
      patterns[635] = 33'b1001100000110110_0_0_00_000_000_000_0_0_00;
      patterns[636] = 33'b1010000000110110_0_1_10_011_110_000_0_x_00;
      patterns[637] = 33'b1010100000110110_1_1_10_011_110_000_0_x_00;
      patterns[638] = 33'b1010100000110110_0_0_00_000_000_000_0_0_00;
      patterns[639] = 33'b1011000000110110_0_1_11_011_110_000_0_x_00;
      patterns[640] = 33'b1011100000110110_1_1_11_011_110_000_0_x_00;
      patterns[641] = 33'b1011100000110110_0_0_00_000_000_000_0_0_00;
      patterns[642] = 33'b0101000000110000_0_1_xx_011_xxx_000_0_1_01;
      patterns[643] = 33'b0101100000110000_1_1_xx_011_xxx_000_0_1_01;
      patterns[644] = 33'b0101100000110000_0_0_00_000_000_000_0_0_00;
      patterns[645] = 33'b0100000000110000_0_0_xx_011_000_xxx_1_x_xx;
      patterns[646] = 33'b0100100000110000_1_0_xx_011_000_xxx_1_x_xx;
      patterns[647] = 33'b0100100000110000_0_0_00_000_000_000_0_0_00;
      patterns[648] = 33'b0000000000111001_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[649] = 33'b0000100000111001_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[650] = 33'b0000100000111001_0_0_00_000_000_000_0_0_00;
      patterns[651] = 33'b1000000000110111_0_1_00_011_111_000_0_x_00;
      patterns[652] = 33'b1000100000110111_1_1_00_011_111_000_0_x_00;
      patterns[653] = 33'b1000100000110111_0_0_00_000_000_000_0_0_00;
      patterns[654] = 33'b1001000000110111_0_1_01_011_111_000_0_x_00;
      patterns[655] = 33'b1001100000110111_1_1_01_011_111_000_0_x_00;
      patterns[656] = 33'b1001100000110111_0_0_00_000_000_000_0_0_00;
      patterns[657] = 33'b1010000000110111_0_1_10_011_111_000_0_x_00;
      patterns[658] = 33'b1010100000110111_1_1_10_011_111_000_0_x_00;
      patterns[659] = 33'b1010100000110111_0_0_00_000_000_000_0_0_00;
      patterns[660] = 33'b1011000000110111_0_1_11_011_111_000_0_x_00;
      patterns[661] = 33'b1011100000110111_1_1_11_011_111_000_0_x_00;
      patterns[662] = 33'b1011100000110111_0_0_00_000_000_000_0_0_00;
      patterns[663] = 33'b0101000000110000_0_1_xx_011_xxx_000_0_1_01;
      patterns[664] = 33'b0101100000110000_1_1_xx_011_xxx_000_0_1_01;
      patterns[665] = 33'b0101100000110000_0_0_00_000_000_000_0_0_00;
      patterns[666] = 33'b0100000000110000_0_0_xx_011_000_xxx_1_x_xx;
      patterns[667] = 33'b0100100000110000_1_0_xx_011_000_xxx_1_x_xx;
      patterns[668] = 33'b0100100000110000_0_0_00_000_000_000_0_0_00;
      patterns[669] = 33'b0000000010101000_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[670] = 33'b0000100010101000_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[671] = 33'b0000100010101000_0_0_00_000_000_000_0_0_00;
      patterns[672] = 33'b1000000001000000_0_1_00_100_000_000_0_x_00;
      patterns[673] = 33'b1000100001000000_1_1_00_100_000_000_0_x_00;
      patterns[674] = 33'b1000100001000000_0_0_00_000_000_000_0_0_00;
      patterns[675] = 33'b1001000001000000_0_1_01_100_000_000_0_x_00;
      patterns[676] = 33'b1001100001000000_1_1_01_100_000_000_0_x_00;
      patterns[677] = 33'b1001100001000000_0_0_00_000_000_000_0_0_00;
      patterns[678] = 33'b1010000001000000_0_1_10_100_000_000_0_x_00;
      patterns[679] = 33'b1010100001000000_1_1_10_100_000_000_0_x_00;
      patterns[680] = 33'b1010100001000000_0_0_00_000_000_000_0_0_00;
      patterns[681] = 33'b1011000001000000_0_1_11_100_000_000_0_x_00;
      patterns[682] = 33'b1011100001000000_1_1_11_100_000_000_0_x_00;
      patterns[683] = 33'b1011100001000000_0_0_00_000_000_000_0_0_00;
      patterns[684] = 33'b0101000001000000_0_1_xx_100_xxx_000_0_1_01;
      patterns[685] = 33'b0101100001000000_1_1_xx_100_xxx_000_0_1_01;
      patterns[686] = 33'b0101100001000000_0_0_00_000_000_000_0_0_00;
      patterns[687] = 33'b0100000001000000_0_0_xx_100_000_xxx_1_x_xx;
      patterns[688] = 33'b0100100001000000_1_0_xx_100_000_xxx_1_x_xx;
      patterns[689] = 33'b0100100001000000_0_0_00_000_000_000_0_0_00;
      patterns[690] = 33'b0000000001100000_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[691] = 33'b0000100001100000_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[692] = 33'b0000100001100000_0_0_00_000_000_000_0_0_00;
      patterns[693] = 33'b1000000001000001_0_1_00_100_001_000_0_x_00;
      patterns[694] = 33'b1000100001000001_1_1_00_100_001_000_0_x_00;
      patterns[695] = 33'b1000100001000001_0_0_00_000_000_000_0_0_00;
      patterns[696] = 33'b1001000001000001_0_1_01_100_001_000_0_x_00;
      patterns[697] = 33'b1001100001000001_1_1_01_100_001_000_0_x_00;
      patterns[698] = 33'b1001100001000001_0_0_00_000_000_000_0_0_00;
      patterns[699] = 33'b1010000001000001_0_1_10_100_001_000_0_x_00;
      patterns[700] = 33'b1010100001000001_1_1_10_100_001_000_0_x_00;
      patterns[701] = 33'b1010100001000001_0_0_00_000_000_000_0_0_00;
      patterns[702] = 33'b1011000001000001_0_1_11_100_001_000_0_x_00;
      patterns[703] = 33'b1011100001000001_1_1_11_100_001_000_0_x_00;
      patterns[704] = 33'b1011100001000001_0_0_00_000_000_000_0_0_00;
      patterns[705] = 33'b0101000001000000_0_1_xx_100_xxx_000_0_1_01;
      patterns[706] = 33'b0101100001000000_1_1_xx_100_xxx_000_0_1_01;
      patterns[707] = 33'b0101100001000000_0_0_00_000_000_000_0_0_00;
      patterns[708] = 33'b0100000001000000_0_0_xx_100_000_xxx_1_x_xx;
      patterns[709] = 33'b0100100001000000_1_0_xx_100_000_xxx_1_x_xx;
      patterns[710] = 33'b0100100001000000_0_0_00_000_000_000_0_0_00;
      patterns[711] = 33'b0000000000010101_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[712] = 33'b0000100000010101_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[713] = 33'b0000100000010101_0_0_00_000_000_000_0_0_00;
      patterns[714] = 33'b1000000001000010_0_1_00_100_010_000_0_x_00;
      patterns[715] = 33'b1000100001000010_1_1_00_100_010_000_0_x_00;
      patterns[716] = 33'b1000100001000010_0_0_00_000_000_000_0_0_00;
      patterns[717] = 33'b1001000001000010_0_1_01_100_010_000_0_x_00;
      patterns[718] = 33'b1001100001000010_1_1_01_100_010_000_0_x_00;
      patterns[719] = 33'b1001100001000010_0_0_00_000_000_000_0_0_00;
      patterns[720] = 33'b1010000001000010_0_1_10_100_010_000_0_x_00;
      patterns[721] = 33'b1010100001000010_1_1_10_100_010_000_0_x_00;
      patterns[722] = 33'b1010100001000010_0_0_00_000_000_000_0_0_00;
      patterns[723] = 33'b1011000001000010_0_1_11_100_010_000_0_x_00;
      patterns[724] = 33'b1011100001000010_1_1_11_100_010_000_0_x_00;
      patterns[725] = 33'b1011100001000010_0_0_00_000_000_000_0_0_00;
      patterns[726] = 33'b0101000001000000_0_1_xx_100_xxx_000_0_1_01;
      patterns[727] = 33'b0101100001000000_1_1_xx_100_xxx_000_0_1_01;
      patterns[728] = 33'b0101100001000000_0_0_00_000_000_000_0_0_00;
      patterns[729] = 33'b0100000001000000_0_0_xx_100_000_xxx_1_x_xx;
      patterns[730] = 33'b0100100001000000_1_0_xx_100_000_xxx_1_x_xx;
      patterns[731] = 33'b0100100001000000_0_0_00_000_000_000_0_0_00;
      patterns[732] = 33'b0000000000111000_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[733] = 33'b0000100000111000_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[734] = 33'b0000100000111000_0_0_00_000_000_000_0_0_00;
      patterns[735] = 33'b1000000001000011_0_1_00_100_011_000_0_x_00;
      patterns[736] = 33'b1000100001000011_1_1_00_100_011_000_0_x_00;
      patterns[737] = 33'b1000100001000011_0_0_00_000_000_000_0_0_00;
      patterns[738] = 33'b1001000001000011_0_1_01_100_011_000_0_x_00;
      patterns[739] = 33'b1001100001000011_1_1_01_100_011_000_0_x_00;
      patterns[740] = 33'b1001100001000011_0_0_00_000_000_000_0_0_00;
      patterns[741] = 33'b1010000001000011_0_1_10_100_011_000_0_x_00;
      patterns[742] = 33'b1010100001000011_1_1_10_100_011_000_0_x_00;
      patterns[743] = 33'b1010100001000011_0_0_00_000_000_000_0_0_00;
      patterns[744] = 33'b1011000001000011_0_1_11_100_011_000_0_x_00;
      patterns[745] = 33'b1011100001000011_1_1_11_100_011_000_0_x_00;
      patterns[746] = 33'b1011100001000011_0_0_00_000_000_000_0_0_00;
      patterns[747] = 33'b0101000001000000_0_1_xx_100_xxx_000_0_1_01;
      patterns[748] = 33'b0101100001000000_1_1_xx_100_xxx_000_0_1_01;
      patterns[749] = 33'b0101100001000000_0_0_00_000_000_000_0_0_00;
      patterns[750] = 33'b0100000001000000_0_0_xx_100_000_xxx_1_x_xx;
      patterns[751] = 33'b0100100001000000_1_0_xx_100_000_xxx_1_x_xx;
      patterns[752] = 33'b0100100001000000_0_0_00_000_000_000_0_0_00;
      patterns[753] = 33'b0000000000100000_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[754] = 33'b0000100000100000_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[755] = 33'b0000100000100000_0_0_00_000_000_000_0_0_00;
      patterns[756] = 33'b1000000001000100_0_1_00_100_100_000_0_x_00;
      patterns[757] = 33'b1000100001000100_1_1_00_100_100_000_0_x_00;
      patterns[758] = 33'b1000100001000100_0_0_00_000_000_000_0_0_00;
      patterns[759] = 33'b1001000001000100_0_1_01_100_100_000_0_x_00;
      patterns[760] = 33'b1001100001000100_1_1_01_100_100_000_0_x_00;
      patterns[761] = 33'b1001100001000100_0_0_00_000_000_000_0_0_00;
      patterns[762] = 33'b1010000001000100_0_1_10_100_100_000_0_x_00;
      patterns[763] = 33'b1010100001000100_1_1_10_100_100_000_0_x_00;
      patterns[764] = 33'b1010100001000100_0_0_00_000_000_000_0_0_00;
      patterns[765] = 33'b1011000001000100_0_1_11_100_100_000_0_x_00;
      patterns[766] = 33'b1011100001000100_1_1_11_100_100_000_0_x_00;
      patterns[767] = 33'b1011100001000100_0_0_00_000_000_000_0_0_00;
      patterns[768] = 33'b0101000001000000_0_1_xx_100_xxx_000_0_1_01;
      patterns[769] = 33'b0101100001000000_1_1_xx_100_xxx_000_0_1_01;
      patterns[770] = 33'b0101100001000000_0_0_00_000_000_000_0_0_00;
      patterns[771] = 33'b0100000001000000_0_0_xx_100_000_xxx_1_x_xx;
      patterns[772] = 33'b0100100001000000_1_0_xx_100_000_xxx_1_x_xx;
      patterns[773] = 33'b0100100001000000_0_0_00_000_000_000_0_0_00;
      patterns[774] = 33'b0000000010111010_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[775] = 33'b0000100010111010_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[776] = 33'b0000100010111010_0_0_00_000_000_000_0_0_00;
      patterns[777] = 33'b1000000001000101_0_1_00_100_101_000_0_x_00;
      patterns[778] = 33'b1000100001000101_1_1_00_100_101_000_0_x_00;
      patterns[779] = 33'b1000100001000101_0_0_00_000_000_000_0_0_00;
      patterns[780] = 33'b1001000001000101_0_1_01_100_101_000_0_x_00;
      patterns[781] = 33'b1001100001000101_1_1_01_100_101_000_0_x_00;
      patterns[782] = 33'b1001100001000101_0_0_00_000_000_000_0_0_00;
      patterns[783] = 33'b1010000001000101_0_1_10_100_101_000_0_x_00;
      patterns[784] = 33'b1010100001000101_1_1_10_100_101_000_0_x_00;
      patterns[785] = 33'b1010100001000101_0_0_00_000_000_000_0_0_00;
      patterns[786] = 33'b1011000001000101_0_1_11_100_101_000_0_x_00;
      patterns[787] = 33'b1011100001000101_1_1_11_100_101_000_0_x_00;
      patterns[788] = 33'b1011100001000101_0_0_00_000_000_000_0_0_00;
      patterns[789] = 33'b0101000001000000_0_1_xx_100_xxx_000_0_1_01;
      patterns[790] = 33'b0101100001000000_1_1_xx_100_xxx_000_0_1_01;
      patterns[791] = 33'b0101100001000000_0_0_00_000_000_000_0_0_00;
      patterns[792] = 33'b0100000001000000_0_0_xx_100_000_xxx_1_x_xx;
      patterns[793] = 33'b0100100001000000_1_0_xx_100_000_xxx_1_x_xx;
      patterns[794] = 33'b0100100001000000_0_0_00_000_000_000_0_0_00;
      patterns[795] = 33'b0000000001110001_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[796] = 33'b0000100001110001_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[797] = 33'b0000100001110001_0_0_00_000_000_000_0_0_00;
      patterns[798] = 33'b1000000001000110_0_1_00_100_110_000_0_x_00;
      patterns[799] = 33'b1000100001000110_1_1_00_100_110_000_0_x_00;
      patterns[800] = 33'b1000100001000110_0_0_00_000_000_000_0_0_00;
      patterns[801] = 33'b1001000001000110_0_1_01_100_110_000_0_x_00;
      patterns[802] = 33'b1001100001000110_1_1_01_100_110_000_0_x_00;
      patterns[803] = 33'b1001100001000110_0_0_00_000_000_000_0_0_00;
      patterns[804] = 33'b1010000001000110_0_1_10_100_110_000_0_x_00;
      patterns[805] = 33'b1010100001000110_1_1_10_100_110_000_0_x_00;
      patterns[806] = 33'b1010100001000110_0_0_00_000_000_000_0_0_00;
      patterns[807] = 33'b1011000001000110_0_1_11_100_110_000_0_x_00;
      patterns[808] = 33'b1011100001000110_1_1_11_100_110_000_0_x_00;
      patterns[809] = 33'b1011100001000110_0_0_00_000_000_000_0_0_00;
      patterns[810] = 33'b0101000001000000_0_1_xx_100_xxx_000_0_1_01;
      patterns[811] = 33'b0101100001000000_1_1_xx_100_xxx_000_0_1_01;
      patterns[812] = 33'b0101100001000000_0_0_00_000_000_000_0_0_00;
      patterns[813] = 33'b0100000001000000_0_0_xx_100_000_xxx_1_x_xx;
      patterns[814] = 33'b0100100001000000_1_0_xx_100_000_xxx_1_x_xx;
      patterns[815] = 33'b0100100001000000_0_0_00_000_000_000_0_0_00;
      patterns[816] = 33'b0000000010011010_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[817] = 33'b0000100010011010_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[818] = 33'b0000100010011010_0_0_00_000_000_000_0_0_00;
      patterns[819] = 33'b1000000001000111_0_1_00_100_111_000_0_x_00;
      patterns[820] = 33'b1000100001000111_1_1_00_100_111_000_0_x_00;
      patterns[821] = 33'b1000100001000111_0_0_00_000_000_000_0_0_00;
      patterns[822] = 33'b1001000001000111_0_1_01_100_111_000_0_x_00;
      patterns[823] = 33'b1001100001000111_1_1_01_100_111_000_0_x_00;
      patterns[824] = 33'b1001100001000111_0_0_00_000_000_000_0_0_00;
      patterns[825] = 33'b1010000001000111_0_1_10_100_111_000_0_x_00;
      patterns[826] = 33'b1010100001000111_1_1_10_100_111_000_0_x_00;
      patterns[827] = 33'b1010100001000111_0_0_00_000_000_000_0_0_00;
      patterns[828] = 33'b1011000001000111_0_1_11_100_111_000_0_x_00;
      patterns[829] = 33'b1011100001000111_1_1_11_100_111_000_0_x_00;
      patterns[830] = 33'b1011100001000111_0_0_00_000_000_000_0_0_00;
      patterns[831] = 33'b0101000001000000_0_1_xx_100_xxx_000_0_1_01;
      patterns[832] = 33'b0101100001000000_1_1_xx_100_xxx_000_0_1_01;
      patterns[833] = 33'b0101100001000000_0_0_00_000_000_000_0_0_00;
      patterns[834] = 33'b0100000001000000_0_0_xx_100_000_xxx_1_x_xx;
      patterns[835] = 33'b0100100001000000_1_0_xx_100_000_xxx_1_x_xx;
      patterns[836] = 33'b0100100001000000_0_0_00_000_000_000_0_0_00;
      patterns[837] = 33'b0000000001010010_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[838] = 33'b0000100001010010_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[839] = 33'b0000100001010010_0_0_00_000_000_000_0_0_00;
      patterns[840] = 33'b1000000001010000_0_1_00_101_000_000_0_x_00;
      patterns[841] = 33'b1000100001010000_1_1_00_101_000_000_0_x_00;
      patterns[842] = 33'b1000100001010000_0_0_00_000_000_000_0_0_00;
      patterns[843] = 33'b1001000001010000_0_1_01_101_000_000_0_x_00;
      patterns[844] = 33'b1001100001010000_1_1_01_101_000_000_0_x_00;
      patterns[845] = 33'b1001100001010000_0_0_00_000_000_000_0_0_00;
      patterns[846] = 33'b1010000001010000_0_1_10_101_000_000_0_x_00;
      patterns[847] = 33'b1010100001010000_1_1_10_101_000_000_0_x_00;
      patterns[848] = 33'b1010100001010000_0_0_00_000_000_000_0_0_00;
      patterns[849] = 33'b1011000001010000_0_1_11_101_000_000_0_x_00;
      patterns[850] = 33'b1011100001010000_1_1_11_101_000_000_0_x_00;
      patterns[851] = 33'b1011100001010000_0_0_00_000_000_000_0_0_00;
      patterns[852] = 33'b0101000001010000_0_1_xx_101_xxx_000_0_1_01;
      patterns[853] = 33'b0101100001010000_1_1_xx_101_xxx_000_0_1_01;
      patterns[854] = 33'b0101100001010000_0_0_00_000_000_000_0_0_00;
      patterns[855] = 33'b0100000001010000_0_0_xx_101_000_xxx_1_x_xx;
      patterns[856] = 33'b0100100001010000_1_0_xx_101_000_xxx_1_x_xx;
      patterns[857] = 33'b0100100001010000_0_0_00_000_000_000_0_0_00;
      patterns[858] = 33'b0000000001111100_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[859] = 33'b0000100001111100_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[860] = 33'b0000100001111100_0_0_00_000_000_000_0_0_00;
      patterns[861] = 33'b1000000001010001_0_1_00_101_001_000_0_x_00;
      patterns[862] = 33'b1000100001010001_1_1_00_101_001_000_0_x_00;
      patterns[863] = 33'b1000100001010001_0_0_00_000_000_000_0_0_00;
      patterns[864] = 33'b1001000001010001_0_1_01_101_001_000_0_x_00;
      patterns[865] = 33'b1001100001010001_1_1_01_101_001_000_0_x_00;
      patterns[866] = 33'b1001100001010001_0_0_00_000_000_000_0_0_00;
      patterns[867] = 33'b1010000001010001_0_1_10_101_001_000_0_x_00;
      patterns[868] = 33'b1010100001010001_1_1_10_101_001_000_0_x_00;
      patterns[869] = 33'b1010100001010001_0_0_00_000_000_000_0_0_00;
      patterns[870] = 33'b1011000001010001_0_1_11_101_001_000_0_x_00;
      patterns[871] = 33'b1011100001010001_1_1_11_101_001_000_0_x_00;
      patterns[872] = 33'b1011100001010001_0_0_00_000_000_000_0_0_00;
      patterns[873] = 33'b0101000001010000_0_1_xx_101_xxx_000_0_1_01;
      patterns[874] = 33'b0101100001010000_1_1_xx_101_xxx_000_0_1_01;
      patterns[875] = 33'b0101100001010000_0_0_00_000_000_000_0_0_00;
      patterns[876] = 33'b0100000001010000_0_0_xx_101_000_xxx_1_x_xx;
      patterns[877] = 33'b0100100001010000_1_0_xx_101_000_xxx_1_x_xx;
      patterns[878] = 33'b0100100001010000_0_0_00_000_000_000_0_0_00;
      patterns[879] = 33'b0000000000101110_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[880] = 33'b0000100000101110_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[881] = 33'b0000100000101110_0_0_00_000_000_000_0_0_00;
      patterns[882] = 33'b1000000001010010_0_1_00_101_010_000_0_x_00;
      patterns[883] = 33'b1000100001010010_1_1_00_101_010_000_0_x_00;
      patterns[884] = 33'b1000100001010010_0_0_00_000_000_000_0_0_00;
      patterns[885] = 33'b1001000001010010_0_1_01_101_010_000_0_x_00;
      patterns[886] = 33'b1001100001010010_1_1_01_101_010_000_0_x_00;
      patterns[887] = 33'b1001100001010010_0_0_00_000_000_000_0_0_00;
      patterns[888] = 33'b1010000001010010_0_1_10_101_010_000_0_x_00;
      patterns[889] = 33'b1010100001010010_1_1_10_101_010_000_0_x_00;
      patterns[890] = 33'b1010100001010010_0_0_00_000_000_000_0_0_00;
      patterns[891] = 33'b1011000001010010_0_1_11_101_010_000_0_x_00;
      patterns[892] = 33'b1011100001010010_1_1_11_101_010_000_0_x_00;
      patterns[893] = 33'b1011100001010010_0_0_00_000_000_000_0_0_00;
      patterns[894] = 33'b0101000001010000_0_1_xx_101_xxx_000_0_1_01;
      patterns[895] = 33'b0101100001010000_1_1_xx_101_xxx_000_0_1_01;
      patterns[896] = 33'b0101100001010000_0_0_00_000_000_000_0_0_00;
      patterns[897] = 33'b0100000001010000_0_0_xx_101_000_xxx_1_x_xx;
      patterns[898] = 33'b0100100001010000_1_0_xx_101_000_xxx_1_x_xx;
      patterns[899] = 33'b0100100001010000_0_0_00_000_000_000_0_0_00;
      patterns[900] = 33'b0000000011000011_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[901] = 33'b0000100011000011_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[902] = 33'b0000100011000011_0_0_00_000_000_000_0_0_00;
      patterns[903] = 33'b1000000001010011_0_1_00_101_011_000_0_x_00;
      patterns[904] = 33'b1000100001010011_1_1_00_101_011_000_0_x_00;
      patterns[905] = 33'b1000100001010011_0_0_00_000_000_000_0_0_00;
      patterns[906] = 33'b1001000001010011_0_1_01_101_011_000_0_x_00;
      patterns[907] = 33'b1001100001010011_1_1_01_101_011_000_0_x_00;
      patterns[908] = 33'b1001100001010011_0_0_00_000_000_000_0_0_00;
      patterns[909] = 33'b1010000001010011_0_1_10_101_011_000_0_x_00;
      patterns[910] = 33'b1010100001010011_1_1_10_101_011_000_0_x_00;
      patterns[911] = 33'b1010100001010011_0_0_00_000_000_000_0_0_00;
      patterns[912] = 33'b1011000001010011_0_1_11_101_011_000_0_x_00;
      patterns[913] = 33'b1011100001010011_1_1_11_101_011_000_0_x_00;
      patterns[914] = 33'b1011100001010011_0_0_00_000_000_000_0_0_00;
      patterns[915] = 33'b0101000001010000_0_1_xx_101_xxx_000_0_1_01;
      patterns[916] = 33'b0101100001010000_1_1_xx_101_xxx_000_0_1_01;
      patterns[917] = 33'b0101100001010000_0_0_00_000_000_000_0_0_00;
      patterns[918] = 33'b0100000001010000_0_0_xx_101_000_xxx_1_x_xx;
      patterns[919] = 33'b0100100001010000_1_0_xx_101_000_xxx_1_x_xx;
      patterns[920] = 33'b0100100001010000_0_0_00_000_000_000_0_0_00;
      patterns[921] = 33'b0000000010010001_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[922] = 33'b0000100010010001_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[923] = 33'b0000100010010001_0_0_00_000_000_000_0_0_00;
      patterns[924] = 33'b1000000001010100_0_1_00_101_100_000_0_x_00;
      patterns[925] = 33'b1000100001010100_1_1_00_101_100_000_0_x_00;
      patterns[926] = 33'b1000100001010100_0_0_00_000_000_000_0_0_00;
      patterns[927] = 33'b1001000001010100_0_1_01_101_100_000_0_x_00;
      patterns[928] = 33'b1001100001010100_1_1_01_101_100_000_0_x_00;
      patterns[929] = 33'b1001100001010100_0_0_00_000_000_000_0_0_00;
      patterns[930] = 33'b1010000001010100_0_1_10_101_100_000_0_x_00;
      patterns[931] = 33'b1010100001010100_1_1_10_101_100_000_0_x_00;
      patterns[932] = 33'b1010100001010100_0_0_00_000_000_000_0_0_00;
      patterns[933] = 33'b1011000001010100_0_1_11_101_100_000_0_x_00;
      patterns[934] = 33'b1011100001010100_1_1_11_101_100_000_0_x_00;
      patterns[935] = 33'b1011100001010100_0_0_00_000_000_000_0_0_00;
      patterns[936] = 33'b0101000001010000_0_1_xx_101_xxx_000_0_1_01;
      patterns[937] = 33'b0101100001010000_1_1_xx_101_xxx_000_0_1_01;
      patterns[938] = 33'b0101100001010000_0_0_00_000_000_000_0_0_00;
      patterns[939] = 33'b0100000001010000_0_0_xx_101_000_xxx_1_x_xx;
      patterns[940] = 33'b0100100001010000_1_0_xx_101_000_xxx_1_x_xx;
      patterns[941] = 33'b0100100001010000_0_0_00_000_000_000_0_0_00;
      patterns[942] = 33'b0000000011010010_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[943] = 33'b0000100011010010_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[944] = 33'b0000100011010010_0_0_00_000_000_000_0_0_00;
      patterns[945] = 33'b1000000001010101_0_1_00_101_101_000_0_x_00;
      patterns[946] = 33'b1000100001010101_1_1_00_101_101_000_0_x_00;
      patterns[947] = 33'b1000100001010101_0_0_00_000_000_000_0_0_00;
      patterns[948] = 33'b1001000001010101_0_1_01_101_101_000_0_x_00;
      patterns[949] = 33'b1001100001010101_1_1_01_101_101_000_0_x_00;
      patterns[950] = 33'b1001100001010101_0_0_00_000_000_000_0_0_00;
      patterns[951] = 33'b1010000001010101_0_1_10_101_101_000_0_x_00;
      patterns[952] = 33'b1010100001010101_1_1_10_101_101_000_0_x_00;
      patterns[953] = 33'b1010100001010101_0_0_00_000_000_000_0_0_00;
      patterns[954] = 33'b1011000001010101_0_1_11_101_101_000_0_x_00;
      patterns[955] = 33'b1011100001010101_1_1_11_101_101_000_0_x_00;
      patterns[956] = 33'b1011100001010101_0_0_00_000_000_000_0_0_00;
      patterns[957] = 33'b0101000001010000_0_1_xx_101_xxx_000_0_1_01;
      patterns[958] = 33'b0101100001010000_1_1_xx_101_xxx_000_0_1_01;
      patterns[959] = 33'b0101100001010000_0_0_00_000_000_000_0_0_00;
      patterns[960] = 33'b0100000001010000_0_0_xx_101_000_xxx_1_x_xx;
      patterns[961] = 33'b0100100001010000_1_0_xx_101_000_xxx_1_x_xx;
      patterns[962] = 33'b0100100001010000_0_0_00_000_000_000_0_0_00;
      patterns[963] = 33'b0000000010110011_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[964] = 33'b0000100010110011_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[965] = 33'b0000100010110011_0_0_00_000_000_000_0_0_00;
      patterns[966] = 33'b1000000001010110_0_1_00_101_110_000_0_x_00;
      patterns[967] = 33'b1000100001010110_1_1_00_101_110_000_0_x_00;
      patterns[968] = 33'b1000100001010110_0_0_00_000_000_000_0_0_00;
      patterns[969] = 33'b1001000001010110_0_1_01_101_110_000_0_x_00;
      patterns[970] = 33'b1001100001010110_1_1_01_101_110_000_0_x_00;
      patterns[971] = 33'b1001100001010110_0_0_00_000_000_000_0_0_00;
      patterns[972] = 33'b1010000001010110_0_1_10_101_110_000_0_x_00;
      patterns[973] = 33'b1010100001010110_1_1_10_101_110_000_0_x_00;
      patterns[974] = 33'b1010100001010110_0_0_00_000_000_000_0_0_00;
      patterns[975] = 33'b1011000001010110_0_1_11_101_110_000_0_x_00;
      patterns[976] = 33'b1011100001010110_1_1_11_101_110_000_0_x_00;
      patterns[977] = 33'b1011100001010110_0_0_00_000_000_000_0_0_00;
      patterns[978] = 33'b0101000001010000_0_1_xx_101_xxx_000_0_1_01;
      patterns[979] = 33'b0101100001010000_1_1_xx_101_xxx_000_0_1_01;
      patterns[980] = 33'b0101100001010000_0_0_00_000_000_000_0_0_00;
      patterns[981] = 33'b0100000001010000_0_0_xx_101_000_xxx_1_x_xx;
      patterns[982] = 33'b0100100001010000_1_0_xx_101_000_xxx_1_x_xx;
      patterns[983] = 33'b0100100001010000_0_0_00_000_000_000_0_0_00;
      patterns[984] = 33'b0000000001010110_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[985] = 33'b0000100001010110_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[986] = 33'b0000100001010110_0_0_00_000_000_000_0_0_00;
      patterns[987] = 33'b1000000001010111_0_1_00_101_111_000_0_x_00;
      patterns[988] = 33'b1000100001010111_1_1_00_101_111_000_0_x_00;
      patterns[989] = 33'b1000100001010111_0_0_00_000_000_000_0_0_00;
      patterns[990] = 33'b1001000001010111_0_1_01_101_111_000_0_x_00;
      patterns[991] = 33'b1001100001010111_1_1_01_101_111_000_0_x_00;
      patterns[992] = 33'b1001100001010111_0_0_00_000_000_000_0_0_00;
      patterns[993] = 33'b1010000001010111_0_1_10_101_111_000_0_x_00;
      patterns[994] = 33'b1010100001010111_1_1_10_101_111_000_0_x_00;
      patterns[995] = 33'b1010100001010111_0_0_00_000_000_000_0_0_00;
      patterns[996] = 33'b1011000001010111_0_1_11_101_111_000_0_x_00;
      patterns[997] = 33'b1011100001010111_1_1_11_101_111_000_0_x_00;
      patterns[998] = 33'b1011100001010111_0_0_00_000_000_000_0_0_00;
      patterns[999] = 33'b0101000001010000_0_1_xx_101_xxx_000_0_1_01;
      patterns[1000] = 33'b0101100001010000_1_1_xx_101_xxx_000_0_1_01;
      patterns[1001] = 33'b0101100001010000_0_0_00_000_000_000_0_0_00;
      patterns[1002] = 33'b0100000001010000_0_0_xx_101_000_xxx_1_x_xx;
      patterns[1003] = 33'b0100100001010000_1_0_xx_101_000_xxx_1_x_xx;
      patterns[1004] = 33'b0100100001010000_0_0_00_000_000_000_0_0_00;
      patterns[1005] = 33'b0000000010101110_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1006] = 33'b0000100010101110_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1007] = 33'b0000100010101110_0_0_00_000_000_000_0_0_00;
      patterns[1008] = 33'b1000000001100000_0_1_00_110_000_000_0_x_00;
      patterns[1009] = 33'b1000100001100000_1_1_00_110_000_000_0_x_00;
      patterns[1010] = 33'b1000100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1011] = 33'b1001000001100000_0_1_01_110_000_000_0_x_00;
      patterns[1012] = 33'b1001100001100000_1_1_01_110_000_000_0_x_00;
      patterns[1013] = 33'b1001100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1014] = 33'b1010000001100000_0_1_10_110_000_000_0_x_00;
      patterns[1015] = 33'b1010100001100000_1_1_10_110_000_000_0_x_00;
      patterns[1016] = 33'b1010100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1017] = 33'b1011000001100000_0_1_11_110_000_000_0_x_00;
      patterns[1018] = 33'b1011100001100000_1_1_11_110_000_000_0_x_00;
      patterns[1019] = 33'b1011100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1020] = 33'b0101000001100000_0_1_xx_110_xxx_000_0_1_01;
      patterns[1021] = 33'b0101100001100000_1_1_xx_110_xxx_000_0_1_01;
      patterns[1022] = 33'b0101100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1023] = 33'b0100000001100000_0_0_xx_110_000_xxx_1_x_xx;
      patterns[1024] = 33'b0100100001100000_1_0_xx_110_000_xxx_1_x_xx;
      patterns[1025] = 33'b0100100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1026] = 33'b0000000010111011_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1027] = 33'b0000100010111011_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1028] = 33'b0000100010111011_0_0_00_000_000_000_0_0_00;
      patterns[1029] = 33'b1000000001100001_0_1_00_110_001_000_0_x_00;
      patterns[1030] = 33'b1000100001100001_1_1_00_110_001_000_0_x_00;
      patterns[1031] = 33'b1000100001100001_0_0_00_000_000_000_0_0_00;
      patterns[1032] = 33'b1001000001100001_0_1_01_110_001_000_0_x_00;
      patterns[1033] = 33'b1001100001100001_1_1_01_110_001_000_0_x_00;
      patterns[1034] = 33'b1001100001100001_0_0_00_000_000_000_0_0_00;
      patterns[1035] = 33'b1010000001100001_0_1_10_110_001_000_0_x_00;
      patterns[1036] = 33'b1010100001100001_1_1_10_110_001_000_0_x_00;
      patterns[1037] = 33'b1010100001100001_0_0_00_000_000_000_0_0_00;
      patterns[1038] = 33'b1011000001100001_0_1_11_110_001_000_0_x_00;
      patterns[1039] = 33'b1011100001100001_1_1_11_110_001_000_0_x_00;
      patterns[1040] = 33'b1011100001100001_0_0_00_000_000_000_0_0_00;
      patterns[1041] = 33'b0101000001100000_0_1_xx_110_xxx_000_0_1_01;
      patterns[1042] = 33'b0101100001100000_1_1_xx_110_xxx_000_0_1_01;
      patterns[1043] = 33'b0101100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1044] = 33'b0100000001100000_0_0_xx_110_000_xxx_1_x_xx;
      patterns[1045] = 33'b0100100001100000_1_0_xx_110_000_xxx_1_x_xx;
      patterns[1046] = 33'b0100100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1047] = 33'b0000000010111001_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1048] = 33'b0000100010111001_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1049] = 33'b0000100010111001_0_0_00_000_000_000_0_0_00;
      patterns[1050] = 33'b1000000001100010_0_1_00_110_010_000_0_x_00;
      patterns[1051] = 33'b1000100001100010_1_1_00_110_010_000_0_x_00;
      patterns[1052] = 33'b1000100001100010_0_0_00_000_000_000_0_0_00;
      patterns[1053] = 33'b1001000001100010_0_1_01_110_010_000_0_x_00;
      patterns[1054] = 33'b1001100001100010_1_1_01_110_010_000_0_x_00;
      patterns[1055] = 33'b1001100001100010_0_0_00_000_000_000_0_0_00;
      patterns[1056] = 33'b1010000001100010_0_1_10_110_010_000_0_x_00;
      patterns[1057] = 33'b1010100001100010_1_1_10_110_010_000_0_x_00;
      patterns[1058] = 33'b1010100001100010_0_0_00_000_000_000_0_0_00;
      patterns[1059] = 33'b1011000001100010_0_1_11_110_010_000_0_x_00;
      patterns[1060] = 33'b1011100001100010_1_1_11_110_010_000_0_x_00;
      patterns[1061] = 33'b1011100001100010_0_0_00_000_000_000_0_0_00;
      patterns[1062] = 33'b0101000001100000_0_1_xx_110_xxx_000_0_1_01;
      patterns[1063] = 33'b0101100001100000_1_1_xx_110_xxx_000_0_1_01;
      patterns[1064] = 33'b0101100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1065] = 33'b0100000001100000_0_0_xx_110_000_xxx_1_x_xx;
      patterns[1066] = 33'b0100100001100000_1_0_xx_110_000_xxx_1_x_xx;
      patterns[1067] = 33'b0100100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1068] = 33'b0000000010000101_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1069] = 33'b0000100010000101_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1070] = 33'b0000100010000101_0_0_00_000_000_000_0_0_00;
      patterns[1071] = 33'b1000000001100011_0_1_00_110_011_000_0_x_00;
      patterns[1072] = 33'b1000100001100011_1_1_00_110_011_000_0_x_00;
      patterns[1073] = 33'b1000100001100011_0_0_00_000_000_000_0_0_00;
      patterns[1074] = 33'b1001000001100011_0_1_01_110_011_000_0_x_00;
      patterns[1075] = 33'b1001100001100011_1_1_01_110_011_000_0_x_00;
      patterns[1076] = 33'b1001100001100011_0_0_00_000_000_000_0_0_00;
      patterns[1077] = 33'b1010000001100011_0_1_10_110_011_000_0_x_00;
      patterns[1078] = 33'b1010100001100011_1_1_10_110_011_000_0_x_00;
      patterns[1079] = 33'b1010100001100011_0_0_00_000_000_000_0_0_00;
      patterns[1080] = 33'b1011000001100011_0_1_11_110_011_000_0_x_00;
      patterns[1081] = 33'b1011100001100011_1_1_11_110_011_000_0_x_00;
      patterns[1082] = 33'b1011100001100011_0_0_00_000_000_000_0_0_00;
      patterns[1083] = 33'b0101000001100000_0_1_xx_110_xxx_000_0_1_01;
      patterns[1084] = 33'b0101100001100000_1_1_xx_110_xxx_000_0_1_01;
      patterns[1085] = 33'b0101100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1086] = 33'b0100000001100000_0_0_xx_110_000_xxx_1_x_xx;
      patterns[1087] = 33'b0100100001100000_1_0_xx_110_000_xxx_1_x_xx;
      patterns[1088] = 33'b0100100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1089] = 33'b0000000011100111_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1090] = 33'b0000100011100111_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1091] = 33'b0000100011100111_0_0_00_000_000_000_0_0_00;
      patterns[1092] = 33'b1000000001100100_0_1_00_110_100_000_0_x_00;
      patterns[1093] = 33'b1000100001100100_1_1_00_110_100_000_0_x_00;
      patterns[1094] = 33'b1000100001100100_0_0_00_000_000_000_0_0_00;
      patterns[1095] = 33'b1001000001100100_0_1_01_110_100_000_0_x_00;
      patterns[1096] = 33'b1001100001100100_1_1_01_110_100_000_0_x_00;
      patterns[1097] = 33'b1001100001100100_0_0_00_000_000_000_0_0_00;
      patterns[1098] = 33'b1010000001100100_0_1_10_110_100_000_0_x_00;
      patterns[1099] = 33'b1010100001100100_1_1_10_110_100_000_0_x_00;
      patterns[1100] = 33'b1010100001100100_0_0_00_000_000_000_0_0_00;
      patterns[1101] = 33'b1011000001100100_0_1_11_110_100_000_0_x_00;
      patterns[1102] = 33'b1011100001100100_1_1_11_110_100_000_0_x_00;
      patterns[1103] = 33'b1011100001100100_0_0_00_000_000_000_0_0_00;
      patterns[1104] = 33'b0101000001100000_0_1_xx_110_xxx_000_0_1_01;
      patterns[1105] = 33'b0101100001100000_1_1_xx_110_xxx_000_0_1_01;
      patterns[1106] = 33'b0101100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1107] = 33'b0100000001100000_0_0_xx_110_000_xxx_1_x_xx;
      patterns[1108] = 33'b0100100001100000_1_0_xx_110_000_xxx_1_x_xx;
      patterns[1109] = 33'b0100100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1110] = 33'b0000000011011011_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1111] = 33'b0000100011011011_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1112] = 33'b0000100011011011_0_0_00_000_000_000_0_0_00;
      patterns[1113] = 33'b1000000001100101_0_1_00_110_101_000_0_x_00;
      patterns[1114] = 33'b1000100001100101_1_1_00_110_101_000_0_x_00;
      patterns[1115] = 33'b1000100001100101_0_0_00_000_000_000_0_0_00;
      patterns[1116] = 33'b1001000001100101_0_1_01_110_101_000_0_x_00;
      patterns[1117] = 33'b1001100001100101_1_1_01_110_101_000_0_x_00;
      patterns[1118] = 33'b1001100001100101_0_0_00_000_000_000_0_0_00;
      patterns[1119] = 33'b1010000001100101_0_1_10_110_101_000_0_x_00;
      patterns[1120] = 33'b1010100001100101_1_1_10_110_101_000_0_x_00;
      patterns[1121] = 33'b1010100001100101_0_0_00_000_000_000_0_0_00;
      patterns[1122] = 33'b1011000001100101_0_1_11_110_101_000_0_x_00;
      patterns[1123] = 33'b1011100001100101_1_1_11_110_101_000_0_x_00;
      patterns[1124] = 33'b1011100001100101_0_0_00_000_000_000_0_0_00;
      patterns[1125] = 33'b0101000001100000_0_1_xx_110_xxx_000_0_1_01;
      patterns[1126] = 33'b0101100001100000_1_1_xx_110_xxx_000_0_1_01;
      patterns[1127] = 33'b0101100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1128] = 33'b0100000001100000_0_0_xx_110_000_xxx_1_x_xx;
      patterns[1129] = 33'b0100100001100000_1_0_xx_110_000_xxx_1_x_xx;
      patterns[1130] = 33'b0100100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1131] = 33'b0000000000111100_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1132] = 33'b0000100000111100_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1133] = 33'b0000100000111100_0_0_00_000_000_000_0_0_00;
      patterns[1134] = 33'b1000000001100110_0_1_00_110_110_000_0_x_00;
      patterns[1135] = 33'b1000100001100110_1_1_00_110_110_000_0_x_00;
      patterns[1136] = 33'b1000100001100110_0_0_00_000_000_000_0_0_00;
      patterns[1137] = 33'b1001000001100110_0_1_01_110_110_000_0_x_00;
      patterns[1138] = 33'b1001100001100110_1_1_01_110_110_000_0_x_00;
      patterns[1139] = 33'b1001100001100110_0_0_00_000_000_000_0_0_00;
      patterns[1140] = 33'b1010000001100110_0_1_10_110_110_000_0_x_00;
      patterns[1141] = 33'b1010100001100110_1_1_10_110_110_000_0_x_00;
      patterns[1142] = 33'b1010100001100110_0_0_00_000_000_000_0_0_00;
      patterns[1143] = 33'b1011000001100110_0_1_11_110_110_000_0_x_00;
      patterns[1144] = 33'b1011100001100110_1_1_11_110_110_000_0_x_00;
      patterns[1145] = 33'b1011100001100110_0_0_00_000_000_000_0_0_00;
      patterns[1146] = 33'b0101000001100000_0_1_xx_110_xxx_000_0_1_01;
      patterns[1147] = 33'b0101100001100000_1_1_xx_110_xxx_000_0_1_01;
      patterns[1148] = 33'b0101100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1149] = 33'b0100000001100000_0_0_xx_110_000_xxx_1_x_xx;
      patterns[1150] = 33'b0100100001100000_1_0_xx_110_000_xxx_1_x_xx;
      patterns[1151] = 33'b0100100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1152] = 33'b0000000010111111_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1153] = 33'b0000100010111111_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1154] = 33'b0000100010111111_0_0_00_000_000_000_0_0_00;
      patterns[1155] = 33'b1000000001100111_0_1_00_110_111_000_0_x_00;
      patterns[1156] = 33'b1000100001100111_1_1_00_110_111_000_0_x_00;
      patterns[1157] = 33'b1000100001100111_0_0_00_000_000_000_0_0_00;
      patterns[1158] = 33'b1001000001100111_0_1_01_110_111_000_0_x_00;
      patterns[1159] = 33'b1001100001100111_1_1_01_110_111_000_0_x_00;
      patterns[1160] = 33'b1001100001100111_0_0_00_000_000_000_0_0_00;
      patterns[1161] = 33'b1010000001100111_0_1_10_110_111_000_0_x_00;
      patterns[1162] = 33'b1010100001100111_1_1_10_110_111_000_0_x_00;
      patterns[1163] = 33'b1010100001100111_0_0_00_000_000_000_0_0_00;
      patterns[1164] = 33'b1011000001100111_0_1_11_110_111_000_0_x_00;
      patterns[1165] = 33'b1011100001100111_1_1_11_110_111_000_0_x_00;
      patterns[1166] = 33'b1011100001100111_0_0_00_000_000_000_0_0_00;
      patterns[1167] = 33'b0101000001100000_0_1_xx_110_xxx_000_0_1_01;
      patterns[1168] = 33'b0101100001100000_1_1_xx_110_xxx_000_0_1_01;
      patterns[1169] = 33'b0101100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1170] = 33'b0100000001100000_0_0_xx_110_000_xxx_1_x_xx;
      patterns[1171] = 33'b0100100001100000_1_0_xx_110_000_xxx_1_x_xx;
      patterns[1172] = 33'b0100100001100000_0_0_00_000_000_000_0_0_00;
      patterns[1173] = 33'b0000000010001000_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1174] = 33'b0000100010001000_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1175] = 33'b0000100010001000_0_0_00_000_000_000_0_0_00;
      patterns[1176] = 33'b1000000001110000_0_1_00_111_000_000_0_x_00;
      patterns[1177] = 33'b1000100001110000_1_1_00_111_000_000_0_x_00;
      patterns[1178] = 33'b1000100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1179] = 33'b1001000001110000_0_1_01_111_000_000_0_x_00;
      patterns[1180] = 33'b1001100001110000_1_1_01_111_000_000_0_x_00;
      patterns[1181] = 33'b1001100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1182] = 33'b1010000001110000_0_1_10_111_000_000_0_x_00;
      patterns[1183] = 33'b1010100001110000_1_1_10_111_000_000_0_x_00;
      patterns[1184] = 33'b1010100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1185] = 33'b1011000001110000_0_1_11_111_000_000_0_x_00;
      patterns[1186] = 33'b1011100001110000_1_1_11_111_000_000_0_x_00;
      patterns[1187] = 33'b1011100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1188] = 33'b0101000001110000_0_1_xx_111_xxx_000_0_1_01;
      patterns[1189] = 33'b0101100001110000_1_1_xx_111_xxx_000_0_1_01;
      patterns[1190] = 33'b0101100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1191] = 33'b0100000001110000_0_0_xx_111_000_xxx_1_x_xx;
      patterns[1192] = 33'b0100100001110000_1_0_xx_111_000_xxx_1_x_xx;
      patterns[1193] = 33'b0100100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1194] = 33'b0000000000000011_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1195] = 33'b0000100000000011_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1196] = 33'b0000100000000011_0_0_00_000_000_000_0_0_00;
      patterns[1197] = 33'b1000000001110001_0_1_00_111_001_000_0_x_00;
      patterns[1198] = 33'b1000100001110001_1_1_00_111_001_000_0_x_00;
      patterns[1199] = 33'b1000100001110001_0_0_00_000_000_000_0_0_00;
      patterns[1200] = 33'b1001000001110001_0_1_01_111_001_000_0_x_00;
      patterns[1201] = 33'b1001100001110001_1_1_01_111_001_000_0_x_00;
      patterns[1202] = 33'b1001100001110001_0_0_00_000_000_000_0_0_00;
      patterns[1203] = 33'b1010000001110001_0_1_10_111_001_000_0_x_00;
      patterns[1204] = 33'b1010100001110001_1_1_10_111_001_000_0_x_00;
      patterns[1205] = 33'b1010100001110001_0_0_00_000_000_000_0_0_00;
      patterns[1206] = 33'b1011000001110001_0_1_11_111_001_000_0_x_00;
      patterns[1207] = 33'b1011100001110001_1_1_11_111_001_000_0_x_00;
      patterns[1208] = 33'b1011100001110001_0_0_00_000_000_000_0_0_00;
      patterns[1209] = 33'b0101000001110000_0_1_xx_111_xxx_000_0_1_01;
      patterns[1210] = 33'b0101100001110000_1_1_xx_111_xxx_000_0_1_01;
      patterns[1211] = 33'b0101100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1212] = 33'b0100000001110000_0_0_xx_111_000_xxx_1_x_xx;
      patterns[1213] = 33'b0100100001110000_1_0_xx_111_000_xxx_1_x_xx;
      patterns[1214] = 33'b0100100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1215] = 33'b0000000011111111_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1216] = 33'b0000100011111111_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1217] = 33'b0000100011111111_0_0_00_000_000_000_0_0_00;
      patterns[1218] = 33'b1000000001110010_0_1_00_111_010_000_0_x_00;
      patterns[1219] = 33'b1000100001110010_1_1_00_111_010_000_0_x_00;
      patterns[1220] = 33'b1000100001110010_0_0_00_000_000_000_0_0_00;
      patterns[1221] = 33'b1001000001110010_0_1_01_111_010_000_0_x_00;
      patterns[1222] = 33'b1001100001110010_1_1_01_111_010_000_0_x_00;
      patterns[1223] = 33'b1001100001110010_0_0_00_000_000_000_0_0_00;
      patterns[1224] = 33'b1010000001110010_0_1_10_111_010_000_0_x_00;
      patterns[1225] = 33'b1010100001110010_1_1_10_111_010_000_0_x_00;
      patterns[1226] = 33'b1010100001110010_0_0_00_000_000_000_0_0_00;
      patterns[1227] = 33'b1011000001110010_0_1_11_111_010_000_0_x_00;
      patterns[1228] = 33'b1011100001110010_1_1_11_111_010_000_0_x_00;
      patterns[1229] = 33'b1011100001110010_0_0_00_000_000_000_0_0_00;
      patterns[1230] = 33'b0101000001110000_0_1_xx_111_xxx_000_0_1_01;
      patterns[1231] = 33'b0101100001110000_1_1_xx_111_xxx_000_0_1_01;
      patterns[1232] = 33'b0101100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1233] = 33'b0100000001110000_0_0_xx_111_000_xxx_1_x_xx;
      patterns[1234] = 33'b0100100001110000_1_0_xx_111_000_xxx_1_x_xx;
      patterns[1235] = 33'b0100100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1236] = 33'b0000000001011010_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1237] = 33'b0000100001011010_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1238] = 33'b0000100001011010_0_0_00_000_000_000_0_0_00;
      patterns[1239] = 33'b1000000001110011_0_1_00_111_011_000_0_x_00;
      patterns[1240] = 33'b1000100001110011_1_1_00_111_011_000_0_x_00;
      patterns[1241] = 33'b1000100001110011_0_0_00_000_000_000_0_0_00;
      patterns[1242] = 33'b1001000001110011_0_1_01_111_011_000_0_x_00;
      patterns[1243] = 33'b1001100001110011_1_1_01_111_011_000_0_x_00;
      patterns[1244] = 33'b1001100001110011_0_0_00_000_000_000_0_0_00;
      patterns[1245] = 33'b1010000001110011_0_1_10_111_011_000_0_x_00;
      patterns[1246] = 33'b1010100001110011_1_1_10_111_011_000_0_x_00;
      patterns[1247] = 33'b1010100001110011_0_0_00_000_000_000_0_0_00;
      patterns[1248] = 33'b1011000001110011_0_1_11_111_011_000_0_x_00;
      patterns[1249] = 33'b1011100001110011_1_1_11_111_011_000_0_x_00;
      patterns[1250] = 33'b1011100001110011_0_0_00_000_000_000_0_0_00;
      patterns[1251] = 33'b0101000001110000_0_1_xx_111_xxx_000_0_1_01;
      patterns[1252] = 33'b0101100001110000_1_1_xx_111_xxx_000_0_1_01;
      patterns[1253] = 33'b0101100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1254] = 33'b0100000001110000_0_0_xx_111_000_xxx_1_x_xx;
      patterns[1255] = 33'b0100100001110000_1_0_xx_111_000_xxx_1_x_xx;
      patterns[1256] = 33'b0100100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1257] = 33'b0000000010010000_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1258] = 33'b0000100010010000_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1259] = 33'b0000100010010000_0_0_00_000_000_000_0_0_00;
      patterns[1260] = 33'b1000000001110100_0_1_00_111_100_000_0_x_00;
      patterns[1261] = 33'b1000100001110100_1_1_00_111_100_000_0_x_00;
      patterns[1262] = 33'b1000100001110100_0_0_00_000_000_000_0_0_00;
      patterns[1263] = 33'b1001000001110100_0_1_01_111_100_000_0_x_00;
      patterns[1264] = 33'b1001100001110100_1_1_01_111_100_000_0_x_00;
      patterns[1265] = 33'b1001100001110100_0_0_00_000_000_000_0_0_00;
      patterns[1266] = 33'b1010000001110100_0_1_10_111_100_000_0_x_00;
      patterns[1267] = 33'b1010100001110100_1_1_10_111_100_000_0_x_00;
      patterns[1268] = 33'b1010100001110100_0_0_00_000_000_000_0_0_00;
      patterns[1269] = 33'b1011000001110100_0_1_11_111_100_000_0_x_00;
      patterns[1270] = 33'b1011100001110100_1_1_11_111_100_000_0_x_00;
      patterns[1271] = 33'b1011100001110100_0_0_00_000_000_000_0_0_00;
      patterns[1272] = 33'b0101000001110000_0_1_xx_111_xxx_000_0_1_01;
      patterns[1273] = 33'b0101100001110000_1_1_xx_111_xxx_000_0_1_01;
      patterns[1274] = 33'b0101100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1275] = 33'b0100000001110000_0_0_xx_111_000_xxx_1_x_xx;
      patterns[1276] = 33'b0100100001110000_1_0_xx_111_000_xxx_1_x_xx;
      patterns[1277] = 33'b0100100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1278] = 33'b0000000001111010_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1279] = 33'b0000100001111010_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1280] = 33'b0000100001111010_0_0_00_000_000_000_0_0_00;
      patterns[1281] = 33'b1000000001110101_0_1_00_111_101_000_0_x_00;
      patterns[1282] = 33'b1000100001110101_1_1_00_111_101_000_0_x_00;
      patterns[1283] = 33'b1000100001110101_0_0_00_000_000_000_0_0_00;
      patterns[1284] = 33'b1001000001110101_0_1_01_111_101_000_0_x_00;
      patterns[1285] = 33'b1001100001110101_1_1_01_111_101_000_0_x_00;
      patterns[1286] = 33'b1001100001110101_0_0_00_000_000_000_0_0_00;
      patterns[1287] = 33'b1010000001110101_0_1_10_111_101_000_0_x_00;
      patterns[1288] = 33'b1010100001110101_1_1_10_111_101_000_0_x_00;
      patterns[1289] = 33'b1010100001110101_0_0_00_000_000_000_0_0_00;
      patterns[1290] = 33'b1011000001110101_0_1_11_111_101_000_0_x_00;
      patterns[1291] = 33'b1011100001110101_1_1_11_111_101_000_0_x_00;
      patterns[1292] = 33'b1011100001110101_0_0_00_000_000_000_0_0_00;
      patterns[1293] = 33'b0101000001110000_0_1_xx_111_xxx_000_0_1_01;
      patterns[1294] = 33'b0101100001110000_1_1_xx_111_xxx_000_0_1_01;
      patterns[1295] = 33'b0101100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1296] = 33'b0100000001110000_0_0_xx_111_000_xxx_1_x_xx;
      patterns[1297] = 33'b0100100001110000_1_0_xx_111_000_xxx_1_x_xx;
      patterns[1298] = 33'b0100100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1299] = 33'b0000000011000100_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1300] = 33'b0000100011000100_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1301] = 33'b0000100011000100_0_0_00_000_000_000_0_0_00;
      patterns[1302] = 33'b1000000001110110_0_1_00_111_110_000_0_x_00;
      patterns[1303] = 33'b1000100001110110_1_1_00_111_110_000_0_x_00;
      patterns[1304] = 33'b1000100001110110_0_0_00_000_000_000_0_0_00;
      patterns[1305] = 33'b1001000001110110_0_1_01_111_110_000_0_x_00;
      patterns[1306] = 33'b1001100001110110_1_1_01_111_110_000_0_x_00;
      patterns[1307] = 33'b1001100001110110_0_0_00_000_000_000_0_0_00;
      patterns[1308] = 33'b1010000001110110_0_1_10_111_110_000_0_x_00;
      patterns[1309] = 33'b1010100001110110_1_1_10_111_110_000_0_x_00;
      patterns[1310] = 33'b1010100001110110_0_0_00_000_000_000_0_0_00;
      patterns[1311] = 33'b1011000001110110_0_1_11_111_110_000_0_x_00;
      patterns[1312] = 33'b1011100001110110_1_1_11_111_110_000_0_x_00;
      patterns[1313] = 33'b1011100001110110_0_0_00_000_000_000_0_0_00;
      patterns[1314] = 33'b0101000001110000_0_1_xx_111_xxx_000_0_1_01;
      patterns[1315] = 33'b0101100001110000_1_1_xx_111_xxx_000_0_1_01;
      patterns[1316] = 33'b0101100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1317] = 33'b0100000001110000_0_0_xx_111_000_xxx_1_x_xx;
      patterns[1318] = 33'b0100100001110000_1_0_xx_111_000_xxx_1_x_xx;
      patterns[1319] = 33'b0100100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1320] = 33'b0000000010101000_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1321] = 33'b0000100010101000_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1322] = 33'b0000100010101000_0_0_00_000_000_000_0_0_00;
      patterns[1323] = 33'b1000000001110111_0_1_00_111_111_000_0_x_00;
      patterns[1324] = 33'b1000100001110111_1_1_00_111_111_000_0_x_00;
      patterns[1325] = 33'b1000100001110111_0_0_00_000_000_000_0_0_00;
      patterns[1326] = 33'b1001000001110111_0_1_01_111_111_000_0_x_00;
      patterns[1327] = 33'b1001100001110111_1_1_01_111_111_000_0_x_00;
      patterns[1328] = 33'b1001100001110111_0_0_00_000_000_000_0_0_00;
      patterns[1329] = 33'b1010000001110111_0_1_10_111_111_000_0_x_00;
      patterns[1330] = 33'b1010100001110111_1_1_10_111_111_000_0_x_00;
      patterns[1331] = 33'b1010100001110111_0_0_00_000_000_000_0_0_00;
      patterns[1332] = 33'b1011000001110111_0_1_11_111_111_000_0_x_00;
      patterns[1333] = 33'b1011100001110111_1_1_11_111_111_000_0_x_00;
      patterns[1334] = 33'b1011100001110111_0_0_00_000_000_000_0_0_00;
      patterns[1335] = 33'b0101000001110000_0_1_xx_111_xxx_000_0_1_01;
      patterns[1336] = 33'b0101100001110000_1_1_xx_111_xxx_000_0_1_01;
      patterns[1337] = 33'b0101100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1338] = 33'b0100000001110000_0_0_xx_111_000_xxx_1_x_xx;
      patterns[1339] = 33'b0100100001110000_1_0_xx_111_000_xxx_1_x_xx;
      patterns[1340] = 33'b0100100001110000_0_0_00_000_000_000_0_0_00;
      patterns[1341] = 33'b0000000001100010_0_1_xx_xxx_xxx_000_0_x_10;
      patterns[1342] = 33'b0000100001100010_1_1_xx_xxx_xxx_000_0_x_10;
      patterns[1343] = 33'b0000100001100010_0_0_00_000_000_000_0_0_00;
      patterns[1344] = 33'b1000000100000000_0_1_00_000_000_001_0_x_00;
      patterns[1345] = 33'b1000100100000000_1_1_00_000_000_001_0_x_00;
      patterns[1346] = 33'b1000100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1347] = 33'b1001000100000000_0_1_01_000_000_001_0_x_00;
      patterns[1348] = 33'b1001100100000000_1_1_01_000_000_001_0_x_00;
      patterns[1349] = 33'b1001100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1350] = 33'b1010000100000000_0_1_10_000_000_001_0_x_00;
      patterns[1351] = 33'b1010100100000000_1_1_10_000_000_001_0_x_00;
      patterns[1352] = 33'b1010100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1353] = 33'b1011000100000000_0_1_11_000_000_001_0_x_00;
      patterns[1354] = 33'b1011100100000000_1_1_11_000_000_001_0_x_00;
      patterns[1355] = 33'b1011100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1356] = 33'b0101000100000000_0_1_xx_000_xxx_001_0_1_01;
      patterns[1357] = 33'b0101100100000000_1_1_xx_000_xxx_001_0_1_01;
      patterns[1358] = 33'b0101100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1359] = 33'b0100000100000000_0_0_xx_000_001_xxx_1_x_xx;
      patterns[1360] = 33'b0100100100000000_1_0_xx_000_001_xxx_1_x_xx;
      patterns[1361] = 33'b0100100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1362] = 33'b0000000110011100_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1363] = 33'b0000100110011100_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1364] = 33'b0000100110011100_0_0_00_000_000_000_0_0_00;
      patterns[1365] = 33'b1000000100000001_0_1_00_000_001_001_0_x_00;
      patterns[1366] = 33'b1000100100000001_1_1_00_000_001_001_0_x_00;
      patterns[1367] = 33'b1000100100000001_0_0_00_000_000_000_0_0_00;
      patterns[1368] = 33'b1001000100000001_0_1_01_000_001_001_0_x_00;
      patterns[1369] = 33'b1001100100000001_1_1_01_000_001_001_0_x_00;
      patterns[1370] = 33'b1001100100000001_0_0_00_000_000_000_0_0_00;
      patterns[1371] = 33'b1010000100000001_0_1_10_000_001_001_0_x_00;
      patterns[1372] = 33'b1010100100000001_1_1_10_000_001_001_0_x_00;
      patterns[1373] = 33'b1010100100000001_0_0_00_000_000_000_0_0_00;
      patterns[1374] = 33'b1011000100000001_0_1_11_000_001_001_0_x_00;
      patterns[1375] = 33'b1011100100000001_1_1_11_000_001_001_0_x_00;
      patterns[1376] = 33'b1011100100000001_0_0_00_000_000_000_0_0_00;
      patterns[1377] = 33'b0101000100000000_0_1_xx_000_xxx_001_0_1_01;
      patterns[1378] = 33'b0101100100000000_1_1_xx_000_xxx_001_0_1_01;
      patterns[1379] = 33'b0101100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1380] = 33'b0100000100000000_0_0_xx_000_001_xxx_1_x_xx;
      patterns[1381] = 33'b0100100100000000_1_0_xx_000_001_xxx_1_x_xx;
      patterns[1382] = 33'b0100100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1383] = 33'b0000000101111111_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1384] = 33'b0000100101111111_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1385] = 33'b0000100101111111_0_0_00_000_000_000_0_0_00;
      patterns[1386] = 33'b1000000100000010_0_1_00_000_010_001_0_x_00;
      patterns[1387] = 33'b1000100100000010_1_1_00_000_010_001_0_x_00;
      patterns[1388] = 33'b1000100100000010_0_0_00_000_000_000_0_0_00;
      patterns[1389] = 33'b1001000100000010_0_1_01_000_010_001_0_x_00;
      patterns[1390] = 33'b1001100100000010_1_1_01_000_010_001_0_x_00;
      patterns[1391] = 33'b1001100100000010_0_0_00_000_000_000_0_0_00;
      patterns[1392] = 33'b1010000100000010_0_1_10_000_010_001_0_x_00;
      patterns[1393] = 33'b1010100100000010_1_1_10_000_010_001_0_x_00;
      patterns[1394] = 33'b1010100100000010_0_0_00_000_000_000_0_0_00;
      patterns[1395] = 33'b1011000100000010_0_1_11_000_010_001_0_x_00;
      patterns[1396] = 33'b1011100100000010_1_1_11_000_010_001_0_x_00;
      patterns[1397] = 33'b1011100100000010_0_0_00_000_000_000_0_0_00;
      patterns[1398] = 33'b0101000100000000_0_1_xx_000_xxx_001_0_1_01;
      patterns[1399] = 33'b0101100100000000_1_1_xx_000_xxx_001_0_1_01;
      patterns[1400] = 33'b0101100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1401] = 33'b0100000100000000_0_0_xx_000_001_xxx_1_x_xx;
      patterns[1402] = 33'b0100100100000000_1_0_xx_000_001_xxx_1_x_xx;
      patterns[1403] = 33'b0100100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1404] = 33'b0000000100110111_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1405] = 33'b0000100100110111_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1406] = 33'b0000100100110111_0_0_00_000_000_000_0_0_00;
      patterns[1407] = 33'b1000000100000011_0_1_00_000_011_001_0_x_00;
      patterns[1408] = 33'b1000100100000011_1_1_00_000_011_001_0_x_00;
      patterns[1409] = 33'b1000100100000011_0_0_00_000_000_000_0_0_00;
      patterns[1410] = 33'b1001000100000011_0_1_01_000_011_001_0_x_00;
      patterns[1411] = 33'b1001100100000011_1_1_01_000_011_001_0_x_00;
      patterns[1412] = 33'b1001100100000011_0_0_00_000_000_000_0_0_00;
      patterns[1413] = 33'b1010000100000011_0_1_10_000_011_001_0_x_00;
      patterns[1414] = 33'b1010100100000011_1_1_10_000_011_001_0_x_00;
      patterns[1415] = 33'b1010100100000011_0_0_00_000_000_000_0_0_00;
      patterns[1416] = 33'b1011000100000011_0_1_11_000_011_001_0_x_00;
      patterns[1417] = 33'b1011100100000011_1_1_11_000_011_001_0_x_00;
      patterns[1418] = 33'b1011100100000011_0_0_00_000_000_000_0_0_00;
      patterns[1419] = 33'b0101000100000000_0_1_xx_000_xxx_001_0_1_01;
      patterns[1420] = 33'b0101100100000000_1_1_xx_000_xxx_001_0_1_01;
      patterns[1421] = 33'b0101100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1422] = 33'b0100000100000000_0_0_xx_000_001_xxx_1_x_xx;
      patterns[1423] = 33'b0100100100000000_1_0_xx_000_001_xxx_1_x_xx;
      patterns[1424] = 33'b0100100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1425] = 33'b0000000101101100_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1426] = 33'b0000100101101100_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1427] = 33'b0000100101101100_0_0_00_000_000_000_0_0_00;
      patterns[1428] = 33'b1000000100000100_0_1_00_000_100_001_0_x_00;
      patterns[1429] = 33'b1000100100000100_1_1_00_000_100_001_0_x_00;
      patterns[1430] = 33'b1000100100000100_0_0_00_000_000_000_0_0_00;
      patterns[1431] = 33'b1001000100000100_0_1_01_000_100_001_0_x_00;
      patterns[1432] = 33'b1001100100000100_1_1_01_000_100_001_0_x_00;
      patterns[1433] = 33'b1001100100000100_0_0_00_000_000_000_0_0_00;
      patterns[1434] = 33'b1010000100000100_0_1_10_000_100_001_0_x_00;
      patterns[1435] = 33'b1010100100000100_1_1_10_000_100_001_0_x_00;
      patterns[1436] = 33'b1010100100000100_0_0_00_000_000_000_0_0_00;
      patterns[1437] = 33'b1011000100000100_0_1_11_000_100_001_0_x_00;
      patterns[1438] = 33'b1011100100000100_1_1_11_000_100_001_0_x_00;
      patterns[1439] = 33'b1011100100000100_0_0_00_000_000_000_0_0_00;
      patterns[1440] = 33'b0101000100000000_0_1_xx_000_xxx_001_0_1_01;
      patterns[1441] = 33'b0101100100000000_1_1_xx_000_xxx_001_0_1_01;
      patterns[1442] = 33'b0101100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1443] = 33'b0100000100000000_0_0_xx_000_001_xxx_1_x_xx;
      patterns[1444] = 33'b0100100100000000_1_0_xx_000_001_xxx_1_x_xx;
      patterns[1445] = 33'b0100100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1446] = 33'b0000000100011011_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1447] = 33'b0000100100011011_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1448] = 33'b0000100100011011_0_0_00_000_000_000_0_0_00;
      patterns[1449] = 33'b1000000100000101_0_1_00_000_101_001_0_x_00;
      patterns[1450] = 33'b1000100100000101_1_1_00_000_101_001_0_x_00;
      patterns[1451] = 33'b1000100100000101_0_0_00_000_000_000_0_0_00;
      patterns[1452] = 33'b1001000100000101_0_1_01_000_101_001_0_x_00;
      patterns[1453] = 33'b1001100100000101_1_1_01_000_101_001_0_x_00;
      patterns[1454] = 33'b1001100100000101_0_0_00_000_000_000_0_0_00;
      patterns[1455] = 33'b1010000100000101_0_1_10_000_101_001_0_x_00;
      patterns[1456] = 33'b1010100100000101_1_1_10_000_101_001_0_x_00;
      patterns[1457] = 33'b1010100100000101_0_0_00_000_000_000_0_0_00;
      patterns[1458] = 33'b1011000100000101_0_1_11_000_101_001_0_x_00;
      patterns[1459] = 33'b1011100100000101_1_1_11_000_101_001_0_x_00;
      patterns[1460] = 33'b1011100100000101_0_0_00_000_000_000_0_0_00;
      patterns[1461] = 33'b0101000100000000_0_1_xx_000_xxx_001_0_1_01;
      patterns[1462] = 33'b0101100100000000_1_1_xx_000_xxx_001_0_1_01;
      patterns[1463] = 33'b0101100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1464] = 33'b0100000100000000_0_0_xx_000_001_xxx_1_x_xx;
      patterns[1465] = 33'b0100100100000000_1_0_xx_000_001_xxx_1_x_xx;
      patterns[1466] = 33'b0100100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1467] = 33'b0000000110001111_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1468] = 33'b0000100110001111_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1469] = 33'b0000100110001111_0_0_00_000_000_000_0_0_00;
      patterns[1470] = 33'b1000000100000110_0_1_00_000_110_001_0_x_00;
      patterns[1471] = 33'b1000100100000110_1_1_00_000_110_001_0_x_00;
      patterns[1472] = 33'b1000100100000110_0_0_00_000_000_000_0_0_00;
      patterns[1473] = 33'b1001000100000110_0_1_01_000_110_001_0_x_00;
      patterns[1474] = 33'b1001100100000110_1_1_01_000_110_001_0_x_00;
      patterns[1475] = 33'b1001100100000110_0_0_00_000_000_000_0_0_00;
      patterns[1476] = 33'b1010000100000110_0_1_10_000_110_001_0_x_00;
      patterns[1477] = 33'b1010100100000110_1_1_10_000_110_001_0_x_00;
      patterns[1478] = 33'b1010100100000110_0_0_00_000_000_000_0_0_00;
      patterns[1479] = 33'b1011000100000110_0_1_11_000_110_001_0_x_00;
      patterns[1480] = 33'b1011100100000110_1_1_11_000_110_001_0_x_00;
      patterns[1481] = 33'b1011100100000110_0_0_00_000_000_000_0_0_00;
      patterns[1482] = 33'b0101000100000000_0_1_xx_000_xxx_001_0_1_01;
      patterns[1483] = 33'b0101100100000000_1_1_xx_000_xxx_001_0_1_01;
      patterns[1484] = 33'b0101100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1485] = 33'b0100000100000000_0_0_xx_000_001_xxx_1_x_xx;
      patterns[1486] = 33'b0100100100000000_1_0_xx_000_001_xxx_1_x_xx;
      patterns[1487] = 33'b0100100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1488] = 33'b0000000101100000_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1489] = 33'b0000100101100000_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1490] = 33'b0000100101100000_0_0_00_000_000_000_0_0_00;
      patterns[1491] = 33'b1000000100000111_0_1_00_000_111_001_0_x_00;
      patterns[1492] = 33'b1000100100000111_1_1_00_000_111_001_0_x_00;
      patterns[1493] = 33'b1000100100000111_0_0_00_000_000_000_0_0_00;
      patterns[1494] = 33'b1001000100000111_0_1_01_000_111_001_0_x_00;
      patterns[1495] = 33'b1001100100000111_1_1_01_000_111_001_0_x_00;
      patterns[1496] = 33'b1001100100000111_0_0_00_000_000_000_0_0_00;
      patterns[1497] = 33'b1010000100000111_0_1_10_000_111_001_0_x_00;
      patterns[1498] = 33'b1010100100000111_1_1_10_000_111_001_0_x_00;
      patterns[1499] = 33'b1010100100000111_0_0_00_000_000_000_0_0_00;
      patterns[1500] = 33'b1011000100000111_0_1_11_000_111_001_0_x_00;
      patterns[1501] = 33'b1011100100000111_1_1_11_000_111_001_0_x_00;
      patterns[1502] = 33'b1011100100000111_0_0_00_000_000_000_0_0_00;
      patterns[1503] = 33'b0101000100000000_0_1_xx_000_xxx_001_0_1_01;
      patterns[1504] = 33'b0101100100000000_1_1_xx_000_xxx_001_0_1_01;
      patterns[1505] = 33'b0101100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1506] = 33'b0100000100000000_0_0_xx_000_001_xxx_1_x_xx;
      patterns[1507] = 33'b0100100100000000_1_0_xx_000_001_xxx_1_x_xx;
      patterns[1508] = 33'b0100100100000000_0_0_00_000_000_000_0_0_00;
      patterns[1509] = 33'b0000000101111111_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1510] = 33'b0000100101111111_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1511] = 33'b0000100101111111_0_0_00_000_000_000_0_0_00;
      patterns[1512] = 33'b1000000100010000_0_1_00_001_000_001_0_x_00;
      patterns[1513] = 33'b1000100100010000_1_1_00_001_000_001_0_x_00;
      patterns[1514] = 33'b1000100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1515] = 33'b1001000100010000_0_1_01_001_000_001_0_x_00;
      patterns[1516] = 33'b1001100100010000_1_1_01_001_000_001_0_x_00;
      patterns[1517] = 33'b1001100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1518] = 33'b1010000100010000_0_1_10_001_000_001_0_x_00;
      patterns[1519] = 33'b1010100100010000_1_1_10_001_000_001_0_x_00;
      patterns[1520] = 33'b1010100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1521] = 33'b1011000100010000_0_1_11_001_000_001_0_x_00;
      patterns[1522] = 33'b1011100100010000_1_1_11_001_000_001_0_x_00;
      patterns[1523] = 33'b1011100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1524] = 33'b0101000100010000_0_1_xx_001_xxx_001_0_1_01;
      patterns[1525] = 33'b0101100100010000_1_1_xx_001_xxx_001_0_1_01;
      patterns[1526] = 33'b0101100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1527] = 33'b0100000100010000_0_0_xx_001_001_xxx_1_x_xx;
      patterns[1528] = 33'b0100100100010000_1_0_xx_001_001_xxx_1_x_xx;
      patterns[1529] = 33'b0100100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1530] = 33'b0000000100101111_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1531] = 33'b0000100100101111_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1532] = 33'b0000100100101111_0_0_00_000_000_000_0_0_00;
      patterns[1533] = 33'b1000000100010001_0_1_00_001_001_001_0_x_00;
      patterns[1534] = 33'b1000100100010001_1_1_00_001_001_001_0_x_00;
      patterns[1535] = 33'b1000100100010001_0_0_00_000_000_000_0_0_00;
      patterns[1536] = 33'b1001000100010001_0_1_01_001_001_001_0_x_00;
      patterns[1537] = 33'b1001100100010001_1_1_01_001_001_001_0_x_00;
      patterns[1538] = 33'b1001100100010001_0_0_00_000_000_000_0_0_00;
      patterns[1539] = 33'b1010000100010001_0_1_10_001_001_001_0_x_00;
      patterns[1540] = 33'b1010100100010001_1_1_10_001_001_001_0_x_00;
      patterns[1541] = 33'b1010100100010001_0_0_00_000_000_000_0_0_00;
      patterns[1542] = 33'b1011000100010001_0_1_11_001_001_001_0_x_00;
      patterns[1543] = 33'b1011100100010001_1_1_11_001_001_001_0_x_00;
      patterns[1544] = 33'b1011100100010001_0_0_00_000_000_000_0_0_00;
      patterns[1545] = 33'b0101000100010000_0_1_xx_001_xxx_001_0_1_01;
      patterns[1546] = 33'b0101100100010000_1_1_xx_001_xxx_001_0_1_01;
      patterns[1547] = 33'b0101100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1548] = 33'b0100000100010000_0_0_xx_001_001_xxx_1_x_xx;
      patterns[1549] = 33'b0100100100010000_1_0_xx_001_001_xxx_1_x_xx;
      patterns[1550] = 33'b0100100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1551] = 33'b0000000100100101_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1552] = 33'b0000100100100101_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1553] = 33'b0000100100100101_0_0_00_000_000_000_0_0_00;
      patterns[1554] = 33'b1000000100010010_0_1_00_001_010_001_0_x_00;
      patterns[1555] = 33'b1000100100010010_1_1_00_001_010_001_0_x_00;
      patterns[1556] = 33'b1000100100010010_0_0_00_000_000_000_0_0_00;
      patterns[1557] = 33'b1001000100010010_0_1_01_001_010_001_0_x_00;
      patterns[1558] = 33'b1001100100010010_1_1_01_001_010_001_0_x_00;
      patterns[1559] = 33'b1001100100010010_0_0_00_000_000_000_0_0_00;
      patterns[1560] = 33'b1010000100010010_0_1_10_001_010_001_0_x_00;
      patterns[1561] = 33'b1010100100010010_1_1_10_001_010_001_0_x_00;
      patterns[1562] = 33'b1010100100010010_0_0_00_000_000_000_0_0_00;
      patterns[1563] = 33'b1011000100010010_0_1_11_001_010_001_0_x_00;
      patterns[1564] = 33'b1011100100010010_1_1_11_001_010_001_0_x_00;
      patterns[1565] = 33'b1011100100010010_0_0_00_000_000_000_0_0_00;
      patterns[1566] = 33'b0101000100010000_0_1_xx_001_xxx_001_0_1_01;
      patterns[1567] = 33'b0101100100010000_1_1_xx_001_xxx_001_0_1_01;
      patterns[1568] = 33'b0101100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1569] = 33'b0100000100010000_0_0_xx_001_001_xxx_1_x_xx;
      patterns[1570] = 33'b0100100100010000_1_0_xx_001_001_xxx_1_x_xx;
      patterns[1571] = 33'b0100100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1572] = 33'b0000000101000010_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1573] = 33'b0000100101000010_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1574] = 33'b0000100101000010_0_0_00_000_000_000_0_0_00;
      patterns[1575] = 33'b1000000100010011_0_1_00_001_011_001_0_x_00;
      patterns[1576] = 33'b1000100100010011_1_1_00_001_011_001_0_x_00;
      patterns[1577] = 33'b1000100100010011_0_0_00_000_000_000_0_0_00;
      patterns[1578] = 33'b1001000100010011_0_1_01_001_011_001_0_x_00;
      patterns[1579] = 33'b1001100100010011_1_1_01_001_011_001_0_x_00;
      patterns[1580] = 33'b1001100100010011_0_0_00_000_000_000_0_0_00;
      patterns[1581] = 33'b1010000100010011_0_1_10_001_011_001_0_x_00;
      patterns[1582] = 33'b1010100100010011_1_1_10_001_011_001_0_x_00;
      patterns[1583] = 33'b1010100100010011_0_0_00_000_000_000_0_0_00;
      patterns[1584] = 33'b1011000100010011_0_1_11_001_011_001_0_x_00;
      patterns[1585] = 33'b1011100100010011_1_1_11_001_011_001_0_x_00;
      patterns[1586] = 33'b1011100100010011_0_0_00_000_000_000_0_0_00;
      patterns[1587] = 33'b0101000100010000_0_1_xx_001_xxx_001_0_1_01;
      patterns[1588] = 33'b0101100100010000_1_1_xx_001_xxx_001_0_1_01;
      patterns[1589] = 33'b0101100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1590] = 33'b0100000100010000_0_0_xx_001_001_xxx_1_x_xx;
      patterns[1591] = 33'b0100100100010000_1_0_xx_001_001_xxx_1_x_xx;
      patterns[1592] = 33'b0100100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1593] = 33'b0000000101111110_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1594] = 33'b0000100101111110_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1595] = 33'b0000100101111110_0_0_00_000_000_000_0_0_00;
      patterns[1596] = 33'b1000000100010100_0_1_00_001_100_001_0_x_00;
      patterns[1597] = 33'b1000100100010100_1_1_00_001_100_001_0_x_00;
      patterns[1598] = 33'b1000100100010100_0_0_00_000_000_000_0_0_00;
      patterns[1599] = 33'b1001000100010100_0_1_01_001_100_001_0_x_00;
      patterns[1600] = 33'b1001100100010100_1_1_01_001_100_001_0_x_00;
      patterns[1601] = 33'b1001100100010100_0_0_00_000_000_000_0_0_00;
      patterns[1602] = 33'b1010000100010100_0_1_10_001_100_001_0_x_00;
      patterns[1603] = 33'b1010100100010100_1_1_10_001_100_001_0_x_00;
      patterns[1604] = 33'b1010100100010100_0_0_00_000_000_000_0_0_00;
      patterns[1605] = 33'b1011000100010100_0_1_11_001_100_001_0_x_00;
      patterns[1606] = 33'b1011100100010100_1_1_11_001_100_001_0_x_00;
      patterns[1607] = 33'b1011100100010100_0_0_00_000_000_000_0_0_00;
      patterns[1608] = 33'b0101000100010000_0_1_xx_001_xxx_001_0_1_01;
      patterns[1609] = 33'b0101100100010000_1_1_xx_001_xxx_001_0_1_01;
      patterns[1610] = 33'b0101100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1611] = 33'b0100000100010000_0_0_xx_001_001_xxx_1_x_xx;
      patterns[1612] = 33'b0100100100010000_1_0_xx_001_001_xxx_1_x_xx;
      patterns[1613] = 33'b0100100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1614] = 33'b0000000101010110_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1615] = 33'b0000100101010110_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1616] = 33'b0000100101010110_0_0_00_000_000_000_0_0_00;
      patterns[1617] = 33'b1000000100010101_0_1_00_001_101_001_0_x_00;
      patterns[1618] = 33'b1000100100010101_1_1_00_001_101_001_0_x_00;
      patterns[1619] = 33'b1000100100010101_0_0_00_000_000_000_0_0_00;
      patterns[1620] = 33'b1001000100010101_0_1_01_001_101_001_0_x_00;
      patterns[1621] = 33'b1001100100010101_1_1_01_001_101_001_0_x_00;
      patterns[1622] = 33'b1001100100010101_0_0_00_000_000_000_0_0_00;
      patterns[1623] = 33'b1010000100010101_0_1_10_001_101_001_0_x_00;
      patterns[1624] = 33'b1010100100010101_1_1_10_001_101_001_0_x_00;
      patterns[1625] = 33'b1010100100010101_0_0_00_000_000_000_0_0_00;
      patterns[1626] = 33'b1011000100010101_0_1_11_001_101_001_0_x_00;
      patterns[1627] = 33'b1011100100010101_1_1_11_001_101_001_0_x_00;
      patterns[1628] = 33'b1011100100010101_0_0_00_000_000_000_0_0_00;
      patterns[1629] = 33'b0101000100010000_0_1_xx_001_xxx_001_0_1_01;
      patterns[1630] = 33'b0101100100010000_1_1_xx_001_xxx_001_0_1_01;
      patterns[1631] = 33'b0101100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1632] = 33'b0100000100010000_0_0_xx_001_001_xxx_1_x_xx;
      patterns[1633] = 33'b0100100100010000_1_0_xx_001_001_xxx_1_x_xx;
      patterns[1634] = 33'b0100100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1635] = 33'b0000000111111000_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1636] = 33'b0000100111111000_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1637] = 33'b0000100111111000_0_0_00_000_000_000_0_0_00;
      patterns[1638] = 33'b1000000100010110_0_1_00_001_110_001_0_x_00;
      patterns[1639] = 33'b1000100100010110_1_1_00_001_110_001_0_x_00;
      patterns[1640] = 33'b1000100100010110_0_0_00_000_000_000_0_0_00;
      patterns[1641] = 33'b1001000100010110_0_1_01_001_110_001_0_x_00;
      patterns[1642] = 33'b1001100100010110_1_1_01_001_110_001_0_x_00;
      patterns[1643] = 33'b1001100100010110_0_0_00_000_000_000_0_0_00;
      patterns[1644] = 33'b1010000100010110_0_1_10_001_110_001_0_x_00;
      patterns[1645] = 33'b1010100100010110_1_1_10_001_110_001_0_x_00;
      patterns[1646] = 33'b1010100100010110_0_0_00_000_000_000_0_0_00;
      patterns[1647] = 33'b1011000100010110_0_1_11_001_110_001_0_x_00;
      patterns[1648] = 33'b1011100100010110_1_1_11_001_110_001_0_x_00;
      patterns[1649] = 33'b1011100100010110_0_0_00_000_000_000_0_0_00;
      patterns[1650] = 33'b0101000100010000_0_1_xx_001_xxx_001_0_1_01;
      patterns[1651] = 33'b0101100100010000_1_1_xx_001_xxx_001_0_1_01;
      patterns[1652] = 33'b0101100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1653] = 33'b0100000100010000_0_0_xx_001_001_xxx_1_x_xx;
      patterns[1654] = 33'b0100100100010000_1_0_xx_001_001_xxx_1_x_xx;
      patterns[1655] = 33'b0100100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1656] = 33'b0000000100000110_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1657] = 33'b0000100100000110_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1658] = 33'b0000100100000110_0_0_00_000_000_000_0_0_00;
      patterns[1659] = 33'b1000000100010111_0_1_00_001_111_001_0_x_00;
      patterns[1660] = 33'b1000100100010111_1_1_00_001_111_001_0_x_00;
      patterns[1661] = 33'b1000100100010111_0_0_00_000_000_000_0_0_00;
      patterns[1662] = 33'b1001000100010111_0_1_01_001_111_001_0_x_00;
      patterns[1663] = 33'b1001100100010111_1_1_01_001_111_001_0_x_00;
      patterns[1664] = 33'b1001100100010111_0_0_00_000_000_000_0_0_00;
      patterns[1665] = 33'b1010000100010111_0_1_10_001_111_001_0_x_00;
      patterns[1666] = 33'b1010100100010111_1_1_10_001_111_001_0_x_00;
      patterns[1667] = 33'b1010100100010111_0_0_00_000_000_000_0_0_00;
      patterns[1668] = 33'b1011000100010111_0_1_11_001_111_001_0_x_00;
      patterns[1669] = 33'b1011100100010111_1_1_11_001_111_001_0_x_00;
      patterns[1670] = 33'b1011100100010111_0_0_00_000_000_000_0_0_00;
      patterns[1671] = 33'b0101000100010000_0_1_xx_001_xxx_001_0_1_01;
      patterns[1672] = 33'b0101100100010000_1_1_xx_001_xxx_001_0_1_01;
      patterns[1673] = 33'b0101100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1674] = 33'b0100000100010000_0_0_xx_001_001_xxx_1_x_xx;
      patterns[1675] = 33'b0100100100010000_1_0_xx_001_001_xxx_1_x_xx;
      patterns[1676] = 33'b0100100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1677] = 33'b0000000111100001_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1678] = 33'b0000100111100001_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1679] = 33'b0000100111100001_0_0_00_000_000_000_0_0_00;
      patterns[1680] = 33'b1000000100100000_0_1_00_010_000_001_0_x_00;
      patterns[1681] = 33'b1000100100100000_1_1_00_010_000_001_0_x_00;
      patterns[1682] = 33'b1000100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1683] = 33'b1001000100100000_0_1_01_010_000_001_0_x_00;
      patterns[1684] = 33'b1001100100100000_1_1_01_010_000_001_0_x_00;
      patterns[1685] = 33'b1001100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1686] = 33'b1010000100100000_0_1_10_010_000_001_0_x_00;
      patterns[1687] = 33'b1010100100100000_1_1_10_010_000_001_0_x_00;
      patterns[1688] = 33'b1010100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1689] = 33'b1011000100100000_0_1_11_010_000_001_0_x_00;
      patterns[1690] = 33'b1011100100100000_1_1_11_010_000_001_0_x_00;
      patterns[1691] = 33'b1011100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1692] = 33'b0101000100100000_0_1_xx_010_xxx_001_0_1_01;
      patterns[1693] = 33'b0101100100100000_1_1_xx_010_xxx_001_0_1_01;
      patterns[1694] = 33'b0101100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1695] = 33'b0100000100100000_0_0_xx_010_001_xxx_1_x_xx;
      patterns[1696] = 33'b0100100100100000_1_0_xx_010_001_xxx_1_x_xx;
      patterns[1697] = 33'b0100100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1698] = 33'b0000000111001110_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1699] = 33'b0000100111001110_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1700] = 33'b0000100111001110_0_0_00_000_000_000_0_0_00;
      patterns[1701] = 33'b1000000100100001_0_1_00_010_001_001_0_x_00;
      patterns[1702] = 33'b1000100100100001_1_1_00_010_001_001_0_x_00;
      patterns[1703] = 33'b1000100100100001_0_0_00_000_000_000_0_0_00;
      patterns[1704] = 33'b1001000100100001_0_1_01_010_001_001_0_x_00;
      patterns[1705] = 33'b1001100100100001_1_1_01_010_001_001_0_x_00;
      patterns[1706] = 33'b1001100100100001_0_0_00_000_000_000_0_0_00;
      patterns[1707] = 33'b1010000100100001_0_1_10_010_001_001_0_x_00;
      patterns[1708] = 33'b1010100100100001_1_1_10_010_001_001_0_x_00;
      patterns[1709] = 33'b1010100100100001_0_0_00_000_000_000_0_0_00;
      patterns[1710] = 33'b1011000100100001_0_1_11_010_001_001_0_x_00;
      patterns[1711] = 33'b1011100100100001_1_1_11_010_001_001_0_x_00;
      patterns[1712] = 33'b1011100100100001_0_0_00_000_000_000_0_0_00;
      patterns[1713] = 33'b0101000100100000_0_1_xx_010_xxx_001_0_1_01;
      patterns[1714] = 33'b0101100100100000_1_1_xx_010_xxx_001_0_1_01;
      patterns[1715] = 33'b0101100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1716] = 33'b0100000100100000_0_0_xx_010_001_xxx_1_x_xx;
      patterns[1717] = 33'b0100100100100000_1_0_xx_010_001_xxx_1_x_xx;
      patterns[1718] = 33'b0100100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1719] = 33'b0000000110000111_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1720] = 33'b0000100110000111_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1721] = 33'b0000100110000111_0_0_00_000_000_000_0_0_00;
      patterns[1722] = 33'b1000000100100010_0_1_00_010_010_001_0_x_00;
      patterns[1723] = 33'b1000100100100010_1_1_00_010_010_001_0_x_00;
      patterns[1724] = 33'b1000100100100010_0_0_00_000_000_000_0_0_00;
      patterns[1725] = 33'b1001000100100010_0_1_01_010_010_001_0_x_00;
      patterns[1726] = 33'b1001100100100010_1_1_01_010_010_001_0_x_00;
      patterns[1727] = 33'b1001100100100010_0_0_00_000_000_000_0_0_00;
      patterns[1728] = 33'b1010000100100010_0_1_10_010_010_001_0_x_00;
      patterns[1729] = 33'b1010100100100010_1_1_10_010_010_001_0_x_00;
      patterns[1730] = 33'b1010100100100010_0_0_00_000_000_000_0_0_00;
      patterns[1731] = 33'b1011000100100010_0_1_11_010_010_001_0_x_00;
      patterns[1732] = 33'b1011100100100010_1_1_11_010_010_001_0_x_00;
      patterns[1733] = 33'b1011100100100010_0_0_00_000_000_000_0_0_00;
      patterns[1734] = 33'b0101000100100000_0_1_xx_010_xxx_001_0_1_01;
      patterns[1735] = 33'b0101100100100000_1_1_xx_010_xxx_001_0_1_01;
      patterns[1736] = 33'b0101100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1737] = 33'b0100000100100000_0_0_xx_010_001_xxx_1_x_xx;
      patterns[1738] = 33'b0100100100100000_1_0_xx_010_001_xxx_1_x_xx;
      patterns[1739] = 33'b0100100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1740] = 33'b0000000100001000_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1741] = 33'b0000100100001000_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1742] = 33'b0000100100001000_0_0_00_000_000_000_0_0_00;
      patterns[1743] = 33'b1000000100100011_0_1_00_010_011_001_0_x_00;
      patterns[1744] = 33'b1000100100100011_1_1_00_010_011_001_0_x_00;
      patterns[1745] = 33'b1000100100100011_0_0_00_000_000_000_0_0_00;
      patterns[1746] = 33'b1001000100100011_0_1_01_010_011_001_0_x_00;
      patterns[1747] = 33'b1001100100100011_1_1_01_010_011_001_0_x_00;
      patterns[1748] = 33'b1001100100100011_0_0_00_000_000_000_0_0_00;
      patterns[1749] = 33'b1010000100100011_0_1_10_010_011_001_0_x_00;
      patterns[1750] = 33'b1010100100100011_1_1_10_010_011_001_0_x_00;
      patterns[1751] = 33'b1010100100100011_0_0_00_000_000_000_0_0_00;
      patterns[1752] = 33'b1011000100100011_0_1_11_010_011_001_0_x_00;
      patterns[1753] = 33'b1011100100100011_1_1_11_010_011_001_0_x_00;
      patterns[1754] = 33'b1011100100100011_0_0_00_000_000_000_0_0_00;
      patterns[1755] = 33'b0101000100100000_0_1_xx_010_xxx_001_0_1_01;
      patterns[1756] = 33'b0101100100100000_1_1_xx_010_xxx_001_0_1_01;
      patterns[1757] = 33'b0101100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1758] = 33'b0100000100100000_0_0_xx_010_001_xxx_1_x_xx;
      patterns[1759] = 33'b0100100100100000_1_0_xx_010_001_xxx_1_x_xx;
      patterns[1760] = 33'b0100100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1761] = 33'b0000000110011010_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1762] = 33'b0000100110011010_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1763] = 33'b0000100110011010_0_0_00_000_000_000_0_0_00;
      patterns[1764] = 33'b1000000100100100_0_1_00_010_100_001_0_x_00;
      patterns[1765] = 33'b1000100100100100_1_1_00_010_100_001_0_x_00;
      patterns[1766] = 33'b1000100100100100_0_0_00_000_000_000_0_0_00;
      patterns[1767] = 33'b1001000100100100_0_1_01_010_100_001_0_x_00;
      patterns[1768] = 33'b1001100100100100_1_1_01_010_100_001_0_x_00;
      patterns[1769] = 33'b1001100100100100_0_0_00_000_000_000_0_0_00;
      patterns[1770] = 33'b1010000100100100_0_1_10_010_100_001_0_x_00;
      patterns[1771] = 33'b1010100100100100_1_1_10_010_100_001_0_x_00;
      patterns[1772] = 33'b1010100100100100_0_0_00_000_000_000_0_0_00;
      patterns[1773] = 33'b1011000100100100_0_1_11_010_100_001_0_x_00;
      patterns[1774] = 33'b1011100100100100_1_1_11_010_100_001_0_x_00;
      patterns[1775] = 33'b1011100100100100_0_0_00_000_000_000_0_0_00;
      patterns[1776] = 33'b0101000100100000_0_1_xx_010_xxx_001_0_1_01;
      patterns[1777] = 33'b0101100100100000_1_1_xx_010_xxx_001_0_1_01;
      patterns[1778] = 33'b0101100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1779] = 33'b0100000100100000_0_0_xx_010_001_xxx_1_x_xx;
      patterns[1780] = 33'b0100100100100000_1_0_xx_010_001_xxx_1_x_xx;
      patterns[1781] = 33'b0100100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1782] = 33'b0000000111100000_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1783] = 33'b0000100111100000_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1784] = 33'b0000100111100000_0_0_00_000_000_000_0_0_00;
      patterns[1785] = 33'b1000000100100101_0_1_00_010_101_001_0_x_00;
      patterns[1786] = 33'b1000100100100101_1_1_00_010_101_001_0_x_00;
      patterns[1787] = 33'b1000100100100101_0_0_00_000_000_000_0_0_00;
      patterns[1788] = 33'b1001000100100101_0_1_01_010_101_001_0_x_00;
      patterns[1789] = 33'b1001100100100101_1_1_01_010_101_001_0_x_00;
      patterns[1790] = 33'b1001100100100101_0_0_00_000_000_000_0_0_00;
      patterns[1791] = 33'b1010000100100101_0_1_10_010_101_001_0_x_00;
      patterns[1792] = 33'b1010100100100101_1_1_10_010_101_001_0_x_00;
      patterns[1793] = 33'b1010100100100101_0_0_00_000_000_000_0_0_00;
      patterns[1794] = 33'b1011000100100101_0_1_11_010_101_001_0_x_00;
      patterns[1795] = 33'b1011100100100101_1_1_11_010_101_001_0_x_00;
      patterns[1796] = 33'b1011100100100101_0_0_00_000_000_000_0_0_00;
      patterns[1797] = 33'b0101000100100000_0_1_xx_010_xxx_001_0_1_01;
      patterns[1798] = 33'b0101100100100000_1_1_xx_010_xxx_001_0_1_01;
      patterns[1799] = 33'b0101100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1800] = 33'b0100000100100000_0_0_xx_010_001_xxx_1_x_xx;
      patterns[1801] = 33'b0100100100100000_1_0_xx_010_001_xxx_1_x_xx;
      patterns[1802] = 33'b0100100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1803] = 33'b0000000100010000_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1804] = 33'b0000100100010000_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1805] = 33'b0000100100010000_0_0_00_000_000_000_0_0_00;
      patterns[1806] = 33'b1000000100100110_0_1_00_010_110_001_0_x_00;
      patterns[1807] = 33'b1000100100100110_1_1_00_010_110_001_0_x_00;
      patterns[1808] = 33'b1000100100100110_0_0_00_000_000_000_0_0_00;
      patterns[1809] = 33'b1001000100100110_0_1_01_010_110_001_0_x_00;
      patterns[1810] = 33'b1001100100100110_1_1_01_010_110_001_0_x_00;
      patterns[1811] = 33'b1001100100100110_0_0_00_000_000_000_0_0_00;
      patterns[1812] = 33'b1010000100100110_0_1_10_010_110_001_0_x_00;
      patterns[1813] = 33'b1010100100100110_1_1_10_010_110_001_0_x_00;
      patterns[1814] = 33'b1010100100100110_0_0_00_000_000_000_0_0_00;
      patterns[1815] = 33'b1011000100100110_0_1_11_010_110_001_0_x_00;
      patterns[1816] = 33'b1011100100100110_1_1_11_010_110_001_0_x_00;
      patterns[1817] = 33'b1011100100100110_0_0_00_000_000_000_0_0_00;
      patterns[1818] = 33'b0101000100100000_0_1_xx_010_xxx_001_0_1_01;
      patterns[1819] = 33'b0101100100100000_1_1_xx_010_xxx_001_0_1_01;
      patterns[1820] = 33'b0101100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1821] = 33'b0100000100100000_0_0_xx_010_001_xxx_1_x_xx;
      patterns[1822] = 33'b0100100100100000_1_0_xx_010_001_xxx_1_x_xx;
      patterns[1823] = 33'b0100100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1824] = 33'b0000000110111001_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1825] = 33'b0000100110111001_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1826] = 33'b0000100110111001_0_0_00_000_000_000_0_0_00;
      patterns[1827] = 33'b1000000100100111_0_1_00_010_111_001_0_x_00;
      patterns[1828] = 33'b1000100100100111_1_1_00_010_111_001_0_x_00;
      patterns[1829] = 33'b1000100100100111_0_0_00_000_000_000_0_0_00;
      patterns[1830] = 33'b1001000100100111_0_1_01_010_111_001_0_x_00;
      patterns[1831] = 33'b1001100100100111_1_1_01_010_111_001_0_x_00;
      patterns[1832] = 33'b1001100100100111_0_0_00_000_000_000_0_0_00;
      patterns[1833] = 33'b1010000100100111_0_1_10_010_111_001_0_x_00;
      patterns[1834] = 33'b1010100100100111_1_1_10_010_111_001_0_x_00;
      patterns[1835] = 33'b1010100100100111_0_0_00_000_000_000_0_0_00;
      patterns[1836] = 33'b1011000100100111_0_1_11_010_111_001_0_x_00;
      patterns[1837] = 33'b1011100100100111_1_1_11_010_111_001_0_x_00;
      patterns[1838] = 33'b1011100100100111_0_0_00_000_000_000_0_0_00;
      patterns[1839] = 33'b0101000100100000_0_1_xx_010_xxx_001_0_1_01;
      patterns[1840] = 33'b0101100100100000_1_1_xx_010_xxx_001_0_1_01;
      patterns[1841] = 33'b0101100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1842] = 33'b0100000100100000_0_0_xx_010_001_xxx_1_x_xx;
      patterns[1843] = 33'b0100100100100000_1_0_xx_010_001_xxx_1_x_xx;
      patterns[1844] = 33'b0100100100100000_0_0_00_000_000_000_0_0_00;
      patterns[1845] = 33'b0000000111001100_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1846] = 33'b0000100111001100_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1847] = 33'b0000100111001100_0_0_00_000_000_000_0_0_00;
      patterns[1848] = 33'b1000000100110000_0_1_00_011_000_001_0_x_00;
      patterns[1849] = 33'b1000100100110000_1_1_00_011_000_001_0_x_00;
      patterns[1850] = 33'b1000100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1851] = 33'b1001000100110000_0_1_01_011_000_001_0_x_00;
      patterns[1852] = 33'b1001100100110000_1_1_01_011_000_001_0_x_00;
      patterns[1853] = 33'b1001100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1854] = 33'b1010000100110000_0_1_10_011_000_001_0_x_00;
      patterns[1855] = 33'b1010100100110000_1_1_10_011_000_001_0_x_00;
      patterns[1856] = 33'b1010100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1857] = 33'b1011000100110000_0_1_11_011_000_001_0_x_00;
      patterns[1858] = 33'b1011100100110000_1_1_11_011_000_001_0_x_00;
      patterns[1859] = 33'b1011100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1860] = 33'b0101000100110000_0_1_xx_011_xxx_001_0_1_01;
      patterns[1861] = 33'b0101100100110000_1_1_xx_011_xxx_001_0_1_01;
      patterns[1862] = 33'b0101100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1863] = 33'b0100000100110000_0_0_xx_011_001_xxx_1_x_xx;
      patterns[1864] = 33'b0100100100110000_1_0_xx_011_001_xxx_1_x_xx;
      patterns[1865] = 33'b0100100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1866] = 33'b0000000100100001_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1867] = 33'b0000100100100001_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1868] = 33'b0000100100100001_0_0_00_000_000_000_0_0_00;
      patterns[1869] = 33'b1000000100110001_0_1_00_011_001_001_0_x_00;
      patterns[1870] = 33'b1000100100110001_1_1_00_011_001_001_0_x_00;
      patterns[1871] = 33'b1000100100110001_0_0_00_000_000_000_0_0_00;
      patterns[1872] = 33'b1001000100110001_0_1_01_011_001_001_0_x_00;
      patterns[1873] = 33'b1001100100110001_1_1_01_011_001_001_0_x_00;
      patterns[1874] = 33'b1001100100110001_0_0_00_000_000_000_0_0_00;
      patterns[1875] = 33'b1010000100110001_0_1_10_011_001_001_0_x_00;
      patterns[1876] = 33'b1010100100110001_1_1_10_011_001_001_0_x_00;
      patterns[1877] = 33'b1010100100110001_0_0_00_000_000_000_0_0_00;
      patterns[1878] = 33'b1011000100110001_0_1_11_011_001_001_0_x_00;
      patterns[1879] = 33'b1011100100110001_1_1_11_011_001_001_0_x_00;
      patterns[1880] = 33'b1011100100110001_0_0_00_000_000_000_0_0_00;
      patterns[1881] = 33'b0101000100110000_0_1_xx_011_xxx_001_0_1_01;
      patterns[1882] = 33'b0101100100110000_1_1_xx_011_xxx_001_0_1_01;
      patterns[1883] = 33'b0101100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1884] = 33'b0100000100110000_0_0_xx_011_001_xxx_1_x_xx;
      patterns[1885] = 33'b0100100100110000_1_0_xx_011_001_xxx_1_x_xx;
      patterns[1886] = 33'b0100100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1887] = 33'b0000000111011010_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1888] = 33'b0000100111011010_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1889] = 33'b0000100111011010_0_0_00_000_000_000_0_0_00;
      patterns[1890] = 33'b1000000100110010_0_1_00_011_010_001_0_x_00;
      patterns[1891] = 33'b1000100100110010_1_1_00_011_010_001_0_x_00;
      patterns[1892] = 33'b1000100100110010_0_0_00_000_000_000_0_0_00;
      patterns[1893] = 33'b1001000100110010_0_1_01_011_010_001_0_x_00;
      patterns[1894] = 33'b1001100100110010_1_1_01_011_010_001_0_x_00;
      patterns[1895] = 33'b1001100100110010_0_0_00_000_000_000_0_0_00;
      patterns[1896] = 33'b1010000100110010_0_1_10_011_010_001_0_x_00;
      patterns[1897] = 33'b1010100100110010_1_1_10_011_010_001_0_x_00;
      patterns[1898] = 33'b1010100100110010_0_0_00_000_000_000_0_0_00;
      patterns[1899] = 33'b1011000100110010_0_1_11_011_010_001_0_x_00;
      patterns[1900] = 33'b1011100100110010_1_1_11_011_010_001_0_x_00;
      patterns[1901] = 33'b1011100100110010_0_0_00_000_000_000_0_0_00;
      patterns[1902] = 33'b0101000100110000_0_1_xx_011_xxx_001_0_1_01;
      patterns[1903] = 33'b0101100100110000_1_1_xx_011_xxx_001_0_1_01;
      patterns[1904] = 33'b0101100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1905] = 33'b0100000100110000_0_0_xx_011_001_xxx_1_x_xx;
      patterns[1906] = 33'b0100100100110000_1_0_xx_011_001_xxx_1_x_xx;
      patterns[1907] = 33'b0100100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1908] = 33'b0000000101010101_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1909] = 33'b0000100101010101_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1910] = 33'b0000100101010101_0_0_00_000_000_000_0_0_00;
      patterns[1911] = 33'b1000000100110011_0_1_00_011_011_001_0_x_00;
      patterns[1912] = 33'b1000100100110011_1_1_00_011_011_001_0_x_00;
      patterns[1913] = 33'b1000100100110011_0_0_00_000_000_000_0_0_00;
      patterns[1914] = 33'b1001000100110011_0_1_01_011_011_001_0_x_00;
      patterns[1915] = 33'b1001100100110011_1_1_01_011_011_001_0_x_00;
      patterns[1916] = 33'b1001100100110011_0_0_00_000_000_000_0_0_00;
      patterns[1917] = 33'b1010000100110011_0_1_10_011_011_001_0_x_00;
      patterns[1918] = 33'b1010100100110011_1_1_10_011_011_001_0_x_00;
      patterns[1919] = 33'b1010100100110011_0_0_00_000_000_000_0_0_00;
      patterns[1920] = 33'b1011000100110011_0_1_11_011_011_001_0_x_00;
      patterns[1921] = 33'b1011100100110011_1_1_11_011_011_001_0_x_00;
      patterns[1922] = 33'b1011100100110011_0_0_00_000_000_000_0_0_00;
      patterns[1923] = 33'b0101000100110000_0_1_xx_011_xxx_001_0_1_01;
      patterns[1924] = 33'b0101100100110000_1_1_xx_011_xxx_001_0_1_01;
      patterns[1925] = 33'b0101100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1926] = 33'b0100000100110000_0_0_xx_011_001_xxx_1_x_xx;
      patterns[1927] = 33'b0100100100110000_1_0_xx_011_001_xxx_1_x_xx;
      patterns[1928] = 33'b0100100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1929] = 33'b0000000111000011_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1930] = 33'b0000100111000011_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1931] = 33'b0000100111000011_0_0_00_000_000_000_0_0_00;
      patterns[1932] = 33'b1000000100110100_0_1_00_011_100_001_0_x_00;
      patterns[1933] = 33'b1000100100110100_1_1_00_011_100_001_0_x_00;
      patterns[1934] = 33'b1000100100110100_0_0_00_000_000_000_0_0_00;
      patterns[1935] = 33'b1001000100110100_0_1_01_011_100_001_0_x_00;
      patterns[1936] = 33'b1001100100110100_1_1_01_011_100_001_0_x_00;
      patterns[1937] = 33'b1001100100110100_0_0_00_000_000_000_0_0_00;
      patterns[1938] = 33'b1010000100110100_0_1_10_011_100_001_0_x_00;
      patterns[1939] = 33'b1010100100110100_1_1_10_011_100_001_0_x_00;
      patterns[1940] = 33'b1010100100110100_0_0_00_000_000_000_0_0_00;
      patterns[1941] = 33'b1011000100110100_0_1_11_011_100_001_0_x_00;
      patterns[1942] = 33'b1011100100110100_1_1_11_011_100_001_0_x_00;
      patterns[1943] = 33'b1011100100110100_0_0_00_000_000_000_0_0_00;
      patterns[1944] = 33'b0101000100110000_0_1_xx_011_xxx_001_0_1_01;
      patterns[1945] = 33'b0101100100110000_1_1_xx_011_xxx_001_0_1_01;
      patterns[1946] = 33'b0101100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1947] = 33'b0100000100110000_0_0_xx_011_001_xxx_1_x_xx;
      patterns[1948] = 33'b0100100100110000_1_0_xx_011_001_xxx_1_x_xx;
      patterns[1949] = 33'b0100100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1950] = 33'b0000000101001011_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1951] = 33'b0000100101001011_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1952] = 33'b0000100101001011_0_0_00_000_000_000_0_0_00;
      patterns[1953] = 33'b1000000100110101_0_1_00_011_101_001_0_x_00;
      patterns[1954] = 33'b1000100100110101_1_1_00_011_101_001_0_x_00;
      patterns[1955] = 33'b1000100100110101_0_0_00_000_000_000_0_0_00;
      patterns[1956] = 33'b1001000100110101_0_1_01_011_101_001_0_x_00;
      patterns[1957] = 33'b1001100100110101_1_1_01_011_101_001_0_x_00;
      patterns[1958] = 33'b1001100100110101_0_0_00_000_000_000_0_0_00;
      patterns[1959] = 33'b1010000100110101_0_1_10_011_101_001_0_x_00;
      patterns[1960] = 33'b1010100100110101_1_1_10_011_101_001_0_x_00;
      patterns[1961] = 33'b1010100100110101_0_0_00_000_000_000_0_0_00;
      patterns[1962] = 33'b1011000100110101_0_1_11_011_101_001_0_x_00;
      patterns[1963] = 33'b1011100100110101_1_1_11_011_101_001_0_x_00;
      patterns[1964] = 33'b1011100100110101_0_0_00_000_000_000_0_0_00;
      patterns[1965] = 33'b0101000100110000_0_1_xx_011_xxx_001_0_1_01;
      patterns[1966] = 33'b0101100100110000_1_1_xx_011_xxx_001_0_1_01;
      patterns[1967] = 33'b0101100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1968] = 33'b0100000100110000_0_0_xx_011_001_xxx_1_x_xx;
      patterns[1969] = 33'b0100100100110000_1_0_xx_011_001_xxx_1_x_xx;
      patterns[1970] = 33'b0100100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1971] = 33'b0000000100011100_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1972] = 33'b0000100100011100_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1973] = 33'b0000100100011100_0_0_00_000_000_000_0_0_00;
      patterns[1974] = 33'b1000000100110110_0_1_00_011_110_001_0_x_00;
      patterns[1975] = 33'b1000100100110110_1_1_00_011_110_001_0_x_00;
      patterns[1976] = 33'b1000100100110110_0_0_00_000_000_000_0_0_00;
      patterns[1977] = 33'b1001000100110110_0_1_01_011_110_001_0_x_00;
      patterns[1978] = 33'b1001100100110110_1_1_01_011_110_001_0_x_00;
      patterns[1979] = 33'b1001100100110110_0_0_00_000_000_000_0_0_00;
      patterns[1980] = 33'b1010000100110110_0_1_10_011_110_001_0_x_00;
      patterns[1981] = 33'b1010100100110110_1_1_10_011_110_001_0_x_00;
      patterns[1982] = 33'b1010100100110110_0_0_00_000_000_000_0_0_00;
      patterns[1983] = 33'b1011000100110110_0_1_11_011_110_001_0_x_00;
      patterns[1984] = 33'b1011100100110110_1_1_11_011_110_001_0_x_00;
      patterns[1985] = 33'b1011100100110110_0_0_00_000_000_000_0_0_00;
      patterns[1986] = 33'b0101000100110000_0_1_xx_011_xxx_001_0_1_01;
      patterns[1987] = 33'b0101100100110000_1_1_xx_011_xxx_001_0_1_01;
      patterns[1988] = 33'b0101100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1989] = 33'b0100000100110000_0_0_xx_011_001_xxx_1_x_xx;
      patterns[1990] = 33'b0100100100110000_1_0_xx_011_001_xxx_1_x_xx;
      patterns[1991] = 33'b0100100100110000_0_0_00_000_000_000_0_0_00;
      patterns[1992] = 33'b0000000101011100_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[1993] = 33'b0000100101011100_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[1994] = 33'b0000100101011100_0_0_00_000_000_000_0_0_00;
      patterns[1995] = 33'b1000000100110111_0_1_00_011_111_001_0_x_00;
      patterns[1996] = 33'b1000100100110111_1_1_00_011_111_001_0_x_00;
      patterns[1997] = 33'b1000100100110111_0_0_00_000_000_000_0_0_00;
      patterns[1998] = 33'b1001000100110111_0_1_01_011_111_001_0_x_00;
      patterns[1999] = 33'b1001100100110111_1_1_01_011_111_001_0_x_00;
      patterns[2000] = 33'b1001100100110111_0_0_00_000_000_000_0_0_00;
      patterns[2001] = 33'b1010000100110111_0_1_10_011_111_001_0_x_00;
      patterns[2002] = 33'b1010100100110111_1_1_10_011_111_001_0_x_00;
      patterns[2003] = 33'b1010100100110111_0_0_00_000_000_000_0_0_00;
      patterns[2004] = 33'b1011000100110111_0_1_11_011_111_001_0_x_00;
      patterns[2005] = 33'b1011100100110111_1_1_11_011_111_001_0_x_00;
      patterns[2006] = 33'b1011100100110111_0_0_00_000_000_000_0_0_00;
      patterns[2007] = 33'b0101000100110000_0_1_xx_011_xxx_001_0_1_01;
      patterns[2008] = 33'b0101100100110000_1_1_xx_011_xxx_001_0_1_01;
      patterns[2009] = 33'b0101100100110000_0_0_00_000_000_000_0_0_00;
      patterns[2010] = 33'b0100000100110000_0_0_xx_011_001_xxx_1_x_xx;
      patterns[2011] = 33'b0100100100110000_1_0_xx_011_001_xxx_1_x_xx;
      patterns[2012] = 33'b0100100100110000_0_0_00_000_000_000_0_0_00;
      patterns[2013] = 33'b0000000111000110_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2014] = 33'b0000100111000110_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2015] = 33'b0000100111000110_0_0_00_000_000_000_0_0_00;
      patterns[2016] = 33'b1000000101000000_0_1_00_100_000_001_0_x_00;
      patterns[2017] = 33'b1000100101000000_1_1_00_100_000_001_0_x_00;
      patterns[2018] = 33'b1000100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2019] = 33'b1001000101000000_0_1_01_100_000_001_0_x_00;
      patterns[2020] = 33'b1001100101000000_1_1_01_100_000_001_0_x_00;
      patterns[2021] = 33'b1001100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2022] = 33'b1010000101000000_0_1_10_100_000_001_0_x_00;
      patterns[2023] = 33'b1010100101000000_1_1_10_100_000_001_0_x_00;
      patterns[2024] = 33'b1010100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2025] = 33'b1011000101000000_0_1_11_100_000_001_0_x_00;
      patterns[2026] = 33'b1011100101000000_1_1_11_100_000_001_0_x_00;
      patterns[2027] = 33'b1011100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2028] = 33'b0101000101000000_0_1_xx_100_xxx_001_0_1_01;
      patterns[2029] = 33'b0101100101000000_1_1_xx_100_xxx_001_0_1_01;
      patterns[2030] = 33'b0101100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2031] = 33'b0100000101000000_0_0_xx_100_001_xxx_1_x_xx;
      patterns[2032] = 33'b0100100101000000_1_0_xx_100_001_xxx_1_x_xx;
      patterns[2033] = 33'b0100100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2034] = 33'b0000000100000100_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2035] = 33'b0000100100000100_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2036] = 33'b0000100100000100_0_0_00_000_000_000_0_0_00;
      patterns[2037] = 33'b1000000101000001_0_1_00_100_001_001_0_x_00;
      patterns[2038] = 33'b1000100101000001_1_1_00_100_001_001_0_x_00;
      patterns[2039] = 33'b1000100101000001_0_0_00_000_000_000_0_0_00;
      patterns[2040] = 33'b1001000101000001_0_1_01_100_001_001_0_x_00;
      patterns[2041] = 33'b1001100101000001_1_1_01_100_001_001_0_x_00;
      patterns[2042] = 33'b1001100101000001_0_0_00_000_000_000_0_0_00;
      patterns[2043] = 33'b1010000101000001_0_1_10_100_001_001_0_x_00;
      patterns[2044] = 33'b1010100101000001_1_1_10_100_001_001_0_x_00;
      patterns[2045] = 33'b1010100101000001_0_0_00_000_000_000_0_0_00;
      patterns[2046] = 33'b1011000101000001_0_1_11_100_001_001_0_x_00;
      patterns[2047] = 33'b1011100101000001_1_1_11_100_001_001_0_x_00;
      patterns[2048] = 33'b1011100101000001_0_0_00_000_000_000_0_0_00;
      patterns[2049] = 33'b0101000101000000_0_1_xx_100_xxx_001_0_1_01;
      patterns[2050] = 33'b0101100101000000_1_1_xx_100_xxx_001_0_1_01;
      patterns[2051] = 33'b0101100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2052] = 33'b0100000101000000_0_0_xx_100_001_xxx_1_x_xx;
      patterns[2053] = 33'b0100100101000000_1_0_xx_100_001_xxx_1_x_xx;
      patterns[2054] = 33'b0100100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2055] = 33'b0000000110000011_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2056] = 33'b0000100110000011_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2057] = 33'b0000100110000011_0_0_00_000_000_000_0_0_00;
      patterns[2058] = 33'b1000000101000010_0_1_00_100_010_001_0_x_00;
      patterns[2059] = 33'b1000100101000010_1_1_00_100_010_001_0_x_00;
      patterns[2060] = 33'b1000100101000010_0_0_00_000_000_000_0_0_00;
      patterns[2061] = 33'b1001000101000010_0_1_01_100_010_001_0_x_00;
      patterns[2062] = 33'b1001100101000010_1_1_01_100_010_001_0_x_00;
      patterns[2063] = 33'b1001100101000010_0_0_00_000_000_000_0_0_00;
      patterns[2064] = 33'b1010000101000010_0_1_10_100_010_001_0_x_00;
      patterns[2065] = 33'b1010100101000010_1_1_10_100_010_001_0_x_00;
      patterns[2066] = 33'b1010100101000010_0_0_00_000_000_000_0_0_00;
      patterns[2067] = 33'b1011000101000010_0_1_11_100_010_001_0_x_00;
      patterns[2068] = 33'b1011100101000010_1_1_11_100_010_001_0_x_00;
      patterns[2069] = 33'b1011100101000010_0_0_00_000_000_000_0_0_00;
      patterns[2070] = 33'b0101000101000000_0_1_xx_100_xxx_001_0_1_01;
      patterns[2071] = 33'b0101100101000000_1_1_xx_100_xxx_001_0_1_01;
      patterns[2072] = 33'b0101100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2073] = 33'b0100000101000000_0_0_xx_100_001_xxx_1_x_xx;
      patterns[2074] = 33'b0100100101000000_1_0_xx_100_001_xxx_1_x_xx;
      patterns[2075] = 33'b0100100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2076] = 33'b0000000110011011_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2077] = 33'b0000100110011011_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2078] = 33'b0000100110011011_0_0_00_000_000_000_0_0_00;
      patterns[2079] = 33'b1000000101000011_0_1_00_100_011_001_0_x_00;
      patterns[2080] = 33'b1000100101000011_1_1_00_100_011_001_0_x_00;
      patterns[2081] = 33'b1000100101000011_0_0_00_000_000_000_0_0_00;
      patterns[2082] = 33'b1001000101000011_0_1_01_100_011_001_0_x_00;
      patterns[2083] = 33'b1001100101000011_1_1_01_100_011_001_0_x_00;
      patterns[2084] = 33'b1001100101000011_0_0_00_000_000_000_0_0_00;
      patterns[2085] = 33'b1010000101000011_0_1_10_100_011_001_0_x_00;
      patterns[2086] = 33'b1010100101000011_1_1_10_100_011_001_0_x_00;
      patterns[2087] = 33'b1010100101000011_0_0_00_000_000_000_0_0_00;
      patterns[2088] = 33'b1011000101000011_0_1_11_100_011_001_0_x_00;
      patterns[2089] = 33'b1011100101000011_1_1_11_100_011_001_0_x_00;
      patterns[2090] = 33'b1011100101000011_0_0_00_000_000_000_0_0_00;
      patterns[2091] = 33'b0101000101000000_0_1_xx_100_xxx_001_0_1_01;
      patterns[2092] = 33'b0101100101000000_1_1_xx_100_xxx_001_0_1_01;
      patterns[2093] = 33'b0101100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2094] = 33'b0100000101000000_0_0_xx_100_001_xxx_1_x_xx;
      patterns[2095] = 33'b0100100101000000_1_0_xx_100_001_xxx_1_x_xx;
      patterns[2096] = 33'b0100100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2097] = 33'b0000000101000111_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2098] = 33'b0000100101000111_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2099] = 33'b0000100101000111_0_0_00_000_000_000_0_0_00;
      patterns[2100] = 33'b1000000101000100_0_1_00_100_100_001_0_x_00;
      patterns[2101] = 33'b1000100101000100_1_1_00_100_100_001_0_x_00;
      patterns[2102] = 33'b1000100101000100_0_0_00_000_000_000_0_0_00;
      patterns[2103] = 33'b1001000101000100_0_1_01_100_100_001_0_x_00;
      patterns[2104] = 33'b1001100101000100_1_1_01_100_100_001_0_x_00;
      patterns[2105] = 33'b1001100101000100_0_0_00_000_000_000_0_0_00;
      patterns[2106] = 33'b1010000101000100_0_1_10_100_100_001_0_x_00;
      patterns[2107] = 33'b1010100101000100_1_1_10_100_100_001_0_x_00;
      patterns[2108] = 33'b1010100101000100_0_0_00_000_000_000_0_0_00;
      patterns[2109] = 33'b1011000101000100_0_1_11_100_100_001_0_x_00;
      patterns[2110] = 33'b1011100101000100_1_1_11_100_100_001_0_x_00;
      patterns[2111] = 33'b1011100101000100_0_0_00_000_000_000_0_0_00;
      patterns[2112] = 33'b0101000101000000_0_1_xx_100_xxx_001_0_1_01;
      patterns[2113] = 33'b0101100101000000_1_1_xx_100_xxx_001_0_1_01;
      patterns[2114] = 33'b0101100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2115] = 33'b0100000101000000_0_0_xx_100_001_xxx_1_x_xx;
      patterns[2116] = 33'b0100100101000000_1_0_xx_100_001_xxx_1_x_xx;
      patterns[2117] = 33'b0100100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2118] = 33'b0000000111011011_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2119] = 33'b0000100111011011_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2120] = 33'b0000100111011011_0_0_00_000_000_000_0_0_00;
      patterns[2121] = 33'b1000000101000101_0_1_00_100_101_001_0_x_00;
      patterns[2122] = 33'b1000100101000101_1_1_00_100_101_001_0_x_00;
      patterns[2123] = 33'b1000100101000101_0_0_00_000_000_000_0_0_00;
      patterns[2124] = 33'b1001000101000101_0_1_01_100_101_001_0_x_00;
      patterns[2125] = 33'b1001100101000101_1_1_01_100_101_001_0_x_00;
      patterns[2126] = 33'b1001100101000101_0_0_00_000_000_000_0_0_00;
      patterns[2127] = 33'b1010000101000101_0_1_10_100_101_001_0_x_00;
      patterns[2128] = 33'b1010100101000101_1_1_10_100_101_001_0_x_00;
      patterns[2129] = 33'b1010100101000101_0_0_00_000_000_000_0_0_00;
      patterns[2130] = 33'b1011000101000101_0_1_11_100_101_001_0_x_00;
      patterns[2131] = 33'b1011100101000101_1_1_11_100_101_001_0_x_00;
      patterns[2132] = 33'b1011100101000101_0_0_00_000_000_000_0_0_00;
      patterns[2133] = 33'b0101000101000000_0_1_xx_100_xxx_001_0_1_01;
      patterns[2134] = 33'b0101100101000000_1_1_xx_100_xxx_001_0_1_01;
      patterns[2135] = 33'b0101100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2136] = 33'b0100000101000000_0_0_xx_100_001_xxx_1_x_xx;
      patterns[2137] = 33'b0100100101000000_1_0_xx_100_001_xxx_1_x_xx;
      patterns[2138] = 33'b0100100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2139] = 33'b0000000100001000_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2140] = 33'b0000100100001000_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2141] = 33'b0000100100001000_0_0_00_000_000_000_0_0_00;
      patterns[2142] = 33'b1000000101000110_0_1_00_100_110_001_0_x_00;
      patterns[2143] = 33'b1000100101000110_1_1_00_100_110_001_0_x_00;
      patterns[2144] = 33'b1000100101000110_0_0_00_000_000_000_0_0_00;
      patterns[2145] = 33'b1001000101000110_0_1_01_100_110_001_0_x_00;
      patterns[2146] = 33'b1001100101000110_1_1_01_100_110_001_0_x_00;
      patterns[2147] = 33'b1001100101000110_0_0_00_000_000_000_0_0_00;
      patterns[2148] = 33'b1010000101000110_0_1_10_100_110_001_0_x_00;
      patterns[2149] = 33'b1010100101000110_1_1_10_100_110_001_0_x_00;
      patterns[2150] = 33'b1010100101000110_0_0_00_000_000_000_0_0_00;
      patterns[2151] = 33'b1011000101000110_0_1_11_100_110_001_0_x_00;
      patterns[2152] = 33'b1011100101000110_1_1_11_100_110_001_0_x_00;
      patterns[2153] = 33'b1011100101000110_0_0_00_000_000_000_0_0_00;
      patterns[2154] = 33'b0101000101000000_0_1_xx_100_xxx_001_0_1_01;
      patterns[2155] = 33'b0101100101000000_1_1_xx_100_xxx_001_0_1_01;
      patterns[2156] = 33'b0101100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2157] = 33'b0100000101000000_0_0_xx_100_001_xxx_1_x_xx;
      patterns[2158] = 33'b0100100101000000_1_0_xx_100_001_xxx_1_x_xx;
      patterns[2159] = 33'b0100100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2160] = 33'b0000000111011111_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2161] = 33'b0000100111011111_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2162] = 33'b0000100111011111_0_0_00_000_000_000_0_0_00;
      patterns[2163] = 33'b1000000101000111_0_1_00_100_111_001_0_x_00;
      patterns[2164] = 33'b1000100101000111_1_1_00_100_111_001_0_x_00;
      patterns[2165] = 33'b1000100101000111_0_0_00_000_000_000_0_0_00;
      patterns[2166] = 33'b1001000101000111_0_1_01_100_111_001_0_x_00;
      patterns[2167] = 33'b1001100101000111_1_1_01_100_111_001_0_x_00;
      patterns[2168] = 33'b1001100101000111_0_0_00_000_000_000_0_0_00;
      patterns[2169] = 33'b1010000101000111_0_1_10_100_111_001_0_x_00;
      patterns[2170] = 33'b1010100101000111_1_1_10_100_111_001_0_x_00;
      patterns[2171] = 33'b1010100101000111_0_0_00_000_000_000_0_0_00;
      patterns[2172] = 33'b1011000101000111_0_1_11_100_111_001_0_x_00;
      patterns[2173] = 33'b1011100101000111_1_1_11_100_111_001_0_x_00;
      patterns[2174] = 33'b1011100101000111_0_0_00_000_000_000_0_0_00;
      patterns[2175] = 33'b0101000101000000_0_1_xx_100_xxx_001_0_1_01;
      patterns[2176] = 33'b0101100101000000_1_1_xx_100_xxx_001_0_1_01;
      patterns[2177] = 33'b0101100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2178] = 33'b0100000101000000_0_0_xx_100_001_xxx_1_x_xx;
      patterns[2179] = 33'b0100100101000000_1_0_xx_100_001_xxx_1_x_xx;
      patterns[2180] = 33'b0100100101000000_0_0_00_000_000_000_0_0_00;
      patterns[2181] = 33'b0000000100100100_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2182] = 33'b0000100100100100_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2183] = 33'b0000100100100100_0_0_00_000_000_000_0_0_00;
      patterns[2184] = 33'b1000000101010000_0_1_00_101_000_001_0_x_00;
      patterns[2185] = 33'b1000100101010000_1_1_00_101_000_001_0_x_00;
      patterns[2186] = 33'b1000100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2187] = 33'b1001000101010000_0_1_01_101_000_001_0_x_00;
      patterns[2188] = 33'b1001100101010000_1_1_01_101_000_001_0_x_00;
      patterns[2189] = 33'b1001100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2190] = 33'b1010000101010000_0_1_10_101_000_001_0_x_00;
      patterns[2191] = 33'b1010100101010000_1_1_10_101_000_001_0_x_00;
      patterns[2192] = 33'b1010100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2193] = 33'b1011000101010000_0_1_11_101_000_001_0_x_00;
      patterns[2194] = 33'b1011100101010000_1_1_11_101_000_001_0_x_00;
      patterns[2195] = 33'b1011100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2196] = 33'b0101000101010000_0_1_xx_101_xxx_001_0_1_01;
      patterns[2197] = 33'b0101100101010000_1_1_xx_101_xxx_001_0_1_01;
      patterns[2198] = 33'b0101100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2199] = 33'b0100000101010000_0_0_xx_101_001_xxx_1_x_xx;
      patterns[2200] = 33'b0100100101010000_1_0_xx_101_001_xxx_1_x_xx;
      patterns[2201] = 33'b0100100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2202] = 33'b0000000100001100_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2203] = 33'b0000100100001100_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2204] = 33'b0000100100001100_0_0_00_000_000_000_0_0_00;
      patterns[2205] = 33'b1000000101010001_0_1_00_101_001_001_0_x_00;
      patterns[2206] = 33'b1000100101010001_1_1_00_101_001_001_0_x_00;
      patterns[2207] = 33'b1000100101010001_0_0_00_000_000_000_0_0_00;
      patterns[2208] = 33'b1001000101010001_0_1_01_101_001_001_0_x_00;
      patterns[2209] = 33'b1001100101010001_1_1_01_101_001_001_0_x_00;
      patterns[2210] = 33'b1001100101010001_0_0_00_000_000_000_0_0_00;
      patterns[2211] = 33'b1010000101010001_0_1_10_101_001_001_0_x_00;
      patterns[2212] = 33'b1010100101010001_1_1_10_101_001_001_0_x_00;
      patterns[2213] = 33'b1010100101010001_0_0_00_000_000_000_0_0_00;
      patterns[2214] = 33'b1011000101010001_0_1_11_101_001_001_0_x_00;
      patterns[2215] = 33'b1011100101010001_1_1_11_101_001_001_0_x_00;
      patterns[2216] = 33'b1011100101010001_0_0_00_000_000_000_0_0_00;
      patterns[2217] = 33'b0101000101010000_0_1_xx_101_xxx_001_0_1_01;
      patterns[2218] = 33'b0101100101010000_1_1_xx_101_xxx_001_0_1_01;
      patterns[2219] = 33'b0101100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2220] = 33'b0100000101010000_0_0_xx_101_001_xxx_1_x_xx;
      patterns[2221] = 33'b0100100101010000_1_0_xx_101_001_xxx_1_x_xx;
      patterns[2222] = 33'b0100100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2223] = 33'b0000000110000000_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2224] = 33'b0000100110000000_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2225] = 33'b0000100110000000_0_0_00_000_000_000_0_0_00;
      patterns[2226] = 33'b1000000101010010_0_1_00_101_010_001_0_x_00;
      patterns[2227] = 33'b1000100101010010_1_1_00_101_010_001_0_x_00;
      patterns[2228] = 33'b1000100101010010_0_0_00_000_000_000_0_0_00;
      patterns[2229] = 33'b1001000101010010_0_1_01_101_010_001_0_x_00;
      patterns[2230] = 33'b1001100101010010_1_1_01_101_010_001_0_x_00;
      patterns[2231] = 33'b1001100101010010_0_0_00_000_000_000_0_0_00;
      patterns[2232] = 33'b1010000101010010_0_1_10_101_010_001_0_x_00;
      patterns[2233] = 33'b1010100101010010_1_1_10_101_010_001_0_x_00;
      patterns[2234] = 33'b1010100101010010_0_0_00_000_000_000_0_0_00;
      patterns[2235] = 33'b1011000101010010_0_1_11_101_010_001_0_x_00;
      patterns[2236] = 33'b1011100101010010_1_1_11_101_010_001_0_x_00;
      patterns[2237] = 33'b1011100101010010_0_0_00_000_000_000_0_0_00;
      patterns[2238] = 33'b0101000101010000_0_1_xx_101_xxx_001_0_1_01;
      patterns[2239] = 33'b0101100101010000_1_1_xx_101_xxx_001_0_1_01;
      patterns[2240] = 33'b0101100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2241] = 33'b0100000101010000_0_0_xx_101_001_xxx_1_x_xx;
      patterns[2242] = 33'b0100100101010000_1_0_xx_101_001_xxx_1_x_xx;
      patterns[2243] = 33'b0100100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2244] = 33'b0000000111110011_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2245] = 33'b0000100111110011_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2246] = 33'b0000100111110011_0_0_00_000_000_000_0_0_00;
      patterns[2247] = 33'b1000000101010011_0_1_00_101_011_001_0_x_00;
      patterns[2248] = 33'b1000100101010011_1_1_00_101_011_001_0_x_00;
      patterns[2249] = 33'b1000100101010011_0_0_00_000_000_000_0_0_00;
      patterns[2250] = 33'b1001000101010011_0_1_01_101_011_001_0_x_00;
      patterns[2251] = 33'b1001100101010011_1_1_01_101_011_001_0_x_00;
      patterns[2252] = 33'b1001100101010011_0_0_00_000_000_000_0_0_00;
      patterns[2253] = 33'b1010000101010011_0_1_10_101_011_001_0_x_00;
      patterns[2254] = 33'b1010100101010011_1_1_10_101_011_001_0_x_00;
      patterns[2255] = 33'b1010100101010011_0_0_00_000_000_000_0_0_00;
      patterns[2256] = 33'b1011000101010011_0_1_11_101_011_001_0_x_00;
      patterns[2257] = 33'b1011100101010011_1_1_11_101_011_001_0_x_00;
      patterns[2258] = 33'b1011100101010011_0_0_00_000_000_000_0_0_00;
      patterns[2259] = 33'b0101000101010000_0_1_xx_101_xxx_001_0_1_01;
      patterns[2260] = 33'b0101100101010000_1_1_xx_101_xxx_001_0_1_01;
      patterns[2261] = 33'b0101100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2262] = 33'b0100000101010000_0_0_xx_101_001_xxx_1_x_xx;
      patterns[2263] = 33'b0100100101010000_1_0_xx_101_001_xxx_1_x_xx;
      patterns[2264] = 33'b0100100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2265] = 33'b0000000111011001_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2266] = 33'b0000100111011001_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2267] = 33'b0000100111011001_0_0_00_000_000_000_0_0_00;
      patterns[2268] = 33'b1000000101010100_0_1_00_101_100_001_0_x_00;
      patterns[2269] = 33'b1000100101010100_1_1_00_101_100_001_0_x_00;
      patterns[2270] = 33'b1000100101010100_0_0_00_000_000_000_0_0_00;
      patterns[2271] = 33'b1001000101010100_0_1_01_101_100_001_0_x_00;
      patterns[2272] = 33'b1001100101010100_1_1_01_101_100_001_0_x_00;
      patterns[2273] = 33'b1001100101010100_0_0_00_000_000_000_0_0_00;
      patterns[2274] = 33'b1010000101010100_0_1_10_101_100_001_0_x_00;
      patterns[2275] = 33'b1010100101010100_1_1_10_101_100_001_0_x_00;
      patterns[2276] = 33'b1010100101010100_0_0_00_000_000_000_0_0_00;
      patterns[2277] = 33'b1011000101010100_0_1_11_101_100_001_0_x_00;
      patterns[2278] = 33'b1011100101010100_1_1_11_101_100_001_0_x_00;
      patterns[2279] = 33'b1011100101010100_0_0_00_000_000_000_0_0_00;
      patterns[2280] = 33'b0101000101010000_0_1_xx_101_xxx_001_0_1_01;
      patterns[2281] = 33'b0101100101010000_1_1_xx_101_xxx_001_0_1_01;
      patterns[2282] = 33'b0101100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2283] = 33'b0100000101010000_0_0_xx_101_001_xxx_1_x_xx;
      patterns[2284] = 33'b0100100101010000_1_0_xx_101_001_xxx_1_x_xx;
      patterns[2285] = 33'b0100100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2286] = 33'b0000000100110101_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2287] = 33'b0000100100110101_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2288] = 33'b0000100100110101_0_0_00_000_000_000_0_0_00;
      patterns[2289] = 33'b1000000101010101_0_1_00_101_101_001_0_x_00;
      patterns[2290] = 33'b1000100101010101_1_1_00_101_101_001_0_x_00;
      patterns[2291] = 33'b1000100101010101_0_0_00_000_000_000_0_0_00;
      patterns[2292] = 33'b1001000101010101_0_1_01_101_101_001_0_x_00;
      patterns[2293] = 33'b1001100101010101_1_1_01_101_101_001_0_x_00;
      patterns[2294] = 33'b1001100101010101_0_0_00_000_000_000_0_0_00;
      patterns[2295] = 33'b1010000101010101_0_1_10_101_101_001_0_x_00;
      patterns[2296] = 33'b1010100101010101_1_1_10_101_101_001_0_x_00;
      patterns[2297] = 33'b1010100101010101_0_0_00_000_000_000_0_0_00;
      patterns[2298] = 33'b1011000101010101_0_1_11_101_101_001_0_x_00;
      patterns[2299] = 33'b1011100101010101_1_1_11_101_101_001_0_x_00;
      patterns[2300] = 33'b1011100101010101_0_0_00_000_000_000_0_0_00;
      patterns[2301] = 33'b0101000101010000_0_1_xx_101_xxx_001_0_1_01;
      patterns[2302] = 33'b0101100101010000_1_1_xx_101_xxx_001_0_1_01;
      patterns[2303] = 33'b0101100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2304] = 33'b0100000101010000_0_0_xx_101_001_xxx_1_x_xx;
      patterns[2305] = 33'b0100100101010000_1_0_xx_101_001_xxx_1_x_xx;
      patterns[2306] = 33'b0100100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2307] = 33'b0000000100100111_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2308] = 33'b0000100100100111_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2309] = 33'b0000100100100111_0_0_00_000_000_000_0_0_00;
      patterns[2310] = 33'b1000000101010110_0_1_00_101_110_001_0_x_00;
      patterns[2311] = 33'b1000100101010110_1_1_00_101_110_001_0_x_00;
      patterns[2312] = 33'b1000100101010110_0_0_00_000_000_000_0_0_00;
      patterns[2313] = 33'b1001000101010110_0_1_01_101_110_001_0_x_00;
      patterns[2314] = 33'b1001100101010110_1_1_01_101_110_001_0_x_00;
      patterns[2315] = 33'b1001100101010110_0_0_00_000_000_000_0_0_00;
      patterns[2316] = 33'b1010000101010110_0_1_10_101_110_001_0_x_00;
      patterns[2317] = 33'b1010100101010110_1_1_10_101_110_001_0_x_00;
      patterns[2318] = 33'b1010100101010110_0_0_00_000_000_000_0_0_00;
      patterns[2319] = 33'b1011000101010110_0_1_11_101_110_001_0_x_00;
      patterns[2320] = 33'b1011100101010110_1_1_11_101_110_001_0_x_00;
      patterns[2321] = 33'b1011100101010110_0_0_00_000_000_000_0_0_00;
      patterns[2322] = 33'b0101000101010000_0_1_xx_101_xxx_001_0_1_01;
      patterns[2323] = 33'b0101100101010000_1_1_xx_101_xxx_001_0_1_01;
      patterns[2324] = 33'b0101100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2325] = 33'b0100000101010000_0_0_xx_101_001_xxx_1_x_xx;
      patterns[2326] = 33'b0100100101010000_1_0_xx_101_001_xxx_1_x_xx;
      patterns[2327] = 33'b0100100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2328] = 33'b0000000101010010_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2329] = 33'b0000100101010010_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2330] = 33'b0000100101010010_0_0_00_000_000_000_0_0_00;
      patterns[2331] = 33'b1000000101010111_0_1_00_101_111_001_0_x_00;
      patterns[2332] = 33'b1000100101010111_1_1_00_101_111_001_0_x_00;
      patterns[2333] = 33'b1000100101010111_0_0_00_000_000_000_0_0_00;
      patterns[2334] = 33'b1001000101010111_0_1_01_101_111_001_0_x_00;
      patterns[2335] = 33'b1001100101010111_1_1_01_101_111_001_0_x_00;
      patterns[2336] = 33'b1001100101010111_0_0_00_000_000_000_0_0_00;
      patterns[2337] = 33'b1010000101010111_0_1_10_101_111_001_0_x_00;
      patterns[2338] = 33'b1010100101010111_1_1_10_101_111_001_0_x_00;
      patterns[2339] = 33'b1010100101010111_0_0_00_000_000_000_0_0_00;
      patterns[2340] = 33'b1011000101010111_0_1_11_101_111_001_0_x_00;
      patterns[2341] = 33'b1011100101010111_1_1_11_101_111_001_0_x_00;
      patterns[2342] = 33'b1011100101010111_0_0_00_000_000_000_0_0_00;
      patterns[2343] = 33'b0101000101010000_0_1_xx_101_xxx_001_0_1_01;
      patterns[2344] = 33'b0101100101010000_1_1_xx_101_xxx_001_0_1_01;
      patterns[2345] = 33'b0101100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2346] = 33'b0100000101010000_0_0_xx_101_001_xxx_1_x_xx;
      patterns[2347] = 33'b0100100101010000_1_0_xx_101_001_xxx_1_x_xx;
      patterns[2348] = 33'b0100100101010000_0_0_00_000_000_000_0_0_00;
      patterns[2349] = 33'b0000000110001010_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2350] = 33'b0000100110001010_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2351] = 33'b0000100110001010_0_0_00_000_000_000_0_0_00;
      patterns[2352] = 33'b1000000101100000_0_1_00_110_000_001_0_x_00;
      patterns[2353] = 33'b1000100101100000_1_1_00_110_000_001_0_x_00;
      patterns[2354] = 33'b1000100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2355] = 33'b1001000101100000_0_1_01_110_000_001_0_x_00;
      patterns[2356] = 33'b1001100101100000_1_1_01_110_000_001_0_x_00;
      patterns[2357] = 33'b1001100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2358] = 33'b1010000101100000_0_1_10_110_000_001_0_x_00;
      patterns[2359] = 33'b1010100101100000_1_1_10_110_000_001_0_x_00;
      patterns[2360] = 33'b1010100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2361] = 33'b1011000101100000_0_1_11_110_000_001_0_x_00;
      patterns[2362] = 33'b1011100101100000_1_1_11_110_000_001_0_x_00;
      patterns[2363] = 33'b1011100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2364] = 33'b0101000101100000_0_1_xx_110_xxx_001_0_1_01;
      patterns[2365] = 33'b0101100101100000_1_1_xx_110_xxx_001_0_1_01;
      patterns[2366] = 33'b0101100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2367] = 33'b0100000101100000_0_0_xx_110_001_xxx_1_x_xx;
      patterns[2368] = 33'b0100100101100000_1_0_xx_110_001_xxx_1_x_xx;
      patterns[2369] = 33'b0100100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2370] = 33'b0000000111010101_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2371] = 33'b0000100111010101_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2372] = 33'b0000100111010101_0_0_00_000_000_000_0_0_00;
      patterns[2373] = 33'b1000000101100001_0_1_00_110_001_001_0_x_00;
      patterns[2374] = 33'b1000100101100001_1_1_00_110_001_001_0_x_00;
      patterns[2375] = 33'b1000100101100001_0_0_00_000_000_000_0_0_00;
      patterns[2376] = 33'b1001000101100001_0_1_01_110_001_001_0_x_00;
      patterns[2377] = 33'b1001100101100001_1_1_01_110_001_001_0_x_00;
      patterns[2378] = 33'b1001100101100001_0_0_00_000_000_000_0_0_00;
      patterns[2379] = 33'b1010000101100001_0_1_10_110_001_001_0_x_00;
      patterns[2380] = 33'b1010100101100001_1_1_10_110_001_001_0_x_00;
      patterns[2381] = 33'b1010100101100001_0_0_00_000_000_000_0_0_00;
      patterns[2382] = 33'b1011000101100001_0_1_11_110_001_001_0_x_00;
      patterns[2383] = 33'b1011100101100001_1_1_11_110_001_001_0_x_00;
      patterns[2384] = 33'b1011100101100001_0_0_00_000_000_000_0_0_00;
      patterns[2385] = 33'b0101000101100000_0_1_xx_110_xxx_001_0_1_01;
      patterns[2386] = 33'b0101100101100000_1_1_xx_110_xxx_001_0_1_01;
      patterns[2387] = 33'b0101100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2388] = 33'b0100000101100000_0_0_xx_110_001_xxx_1_x_xx;
      patterns[2389] = 33'b0100100101100000_1_0_xx_110_001_xxx_1_x_xx;
      patterns[2390] = 33'b0100100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2391] = 33'b0000000100011011_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2392] = 33'b0000100100011011_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2393] = 33'b0000100100011011_0_0_00_000_000_000_0_0_00;
      patterns[2394] = 33'b1000000101100010_0_1_00_110_010_001_0_x_00;
      patterns[2395] = 33'b1000100101100010_1_1_00_110_010_001_0_x_00;
      patterns[2396] = 33'b1000100101100010_0_0_00_000_000_000_0_0_00;
      patterns[2397] = 33'b1001000101100010_0_1_01_110_010_001_0_x_00;
      patterns[2398] = 33'b1001100101100010_1_1_01_110_010_001_0_x_00;
      patterns[2399] = 33'b1001100101100010_0_0_00_000_000_000_0_0_00;
      patterns[2400] = 33'b1010000101100010_0_1_10_110_010_001_0_x_00;
      patterns[2401] = 33'b1010100101100010_1_1_10_110_010_001_0_x_00;
      patterns[2402] = 33'b1010100101100010_0_0_00_000_000_000_0_0_00;
      patterns[2403] = 33'b1011000101100010_0_1_11_110_010_001_0_x_00;
      patterns[2404] = 33'b1011100101100010_1_1_11_110_010_001_0_x_00;
      patterns[2405] = 33'b1011100101100010_0_0_00_000_000_000_0_0_00;
      patterns[2406] = 33'b0101000101100000_0_1_xx_110_xxx_001_0_1_01;
      patterns[2407] = 33'b0101100101100000_1_1_xx_110_xxx_001_0_1_01;
      patterns[2408] = 33'b0101100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2409] = 33'b0100000101100000_0_0_xx_110_001_xxx_1_x_xx;
      patterns[2410] = 33'b0100100101100000_1_0_xx_110_001_xxx_1_x_xx;
      patterns[2411] = 33'b0100100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2412] = 33'b0000000100011010_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2413] = 33'b0000100100011010_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2414] = 33'b0000100100011010_0_0_00_000_000_000_0_0_00;
      patterns[2415] = 33'b1000000101100011_0_1_00_110_011_001_0_x_00;
      patterns[2416] = 33'b1000100101100011_1_1_00_110_011_001_0_x_00;
      patterns[2417] = 33'b1000100101100011_0_0_00_000_000_000_0_0_00;
      patterns[2418] = 33'b1001000101100011_0_1_01_110_011_001_0_x_00;
      patterns[2419] = 33'b1001100101100011_1_1_01_110_011_001_0_x_00;
      patterns[2420] = 33'b1001100101100011_0_0_00_000_000_000_0_0_00;
      patterns[2421] = 33'b1010000101100011_0_1_10_110_011_001_0_x_00;
      patterns[2422] = 33'b1010100101100011_1_1_10_110_011_001_0_x_00;
      patterns[2423] = 33'b1010100101100011_0_0_00_000_000_000_0_0_00;
      patterns[2424] = 33'b1011000101100011_0_1_11_110_011_001_0_x_00;
      patterns[2425] = 33'b1011100101100011_1_1_11_110_011_001_0_x_00;
      patterns[2426] = 33'b1011100101100011_0_0_00_000_000_000_0_0_00;
      patterns[2427] = 33'b0101000101100000_0_1_xx_110_xxx_001_0_1_01;
      patterns[2428] = 33'b0101100101100000_1_1_xx_110_xxx_001_0_1_01;
      patterns[2429] = 33'b0101100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2430] = 33'b0100000101100000_0_0_xx_110_001_xxx_1_x_xx;
      patterns[2431] = 33'b0100100101100000_1_0_xx_110_001_xxx_1_x_xx;
      patterns[2432] = 33'b0100100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2433] = 33'b0000000100100101_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2434] = 33'b0000100100100101_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2435] = 33'b0000100100100101_0_0_00_000_000_000_0_0_00;
      patterns[2436] = 33'b1000000101100100_0_1_00_110_100_001_0_x_00;
      patterns[2437] = 33'b1000100101100100_1_1_00_110_100_001_0_x_00;
      patterns[2438] = 33'b1000100101100100_0_0_00_000_000_000_0_0_00;
      patterns[2439] = 33'b1001000101100100_0_1_01_110_100_001_0_x_00;
      patterns[2440] = 33'b1001100101100100_1_1_01_110_100_001_0_x_00;
      patterns[2441] = 33'b1001100101100100_0_0_00_000_000_000_0_0_00;
      patterns[2442] = 33'b1010000101100100_0_1_10_110_100_001_0_x_00;
      patterns[2443] = 33'b1010100101100100_1_1_10_110_100_001_0_x_00;
      patterns[2444] = 33'b1010100101100100_0_0_00_000_000_000_0_0_00;
      patterns[2445] = 33'b1011000101100100_0_1_11_110_100_001_0_x_00;
      patterns[2446] = 33'b1011100101100100_1_1_11_110_100_001_0_x_00;
      patterns[2447] = 33'b1011100101100100_0_0_00_000_000_000_0_0_00;
      patterns[2448] = 33'b0101000101100000_0_1_xx_110_xxx_001_0_1_01;
      patterns[2449] = 33'b0101100101100000_1_1_xx_110_xxx_001_0_1_01;
      patterns[2450] = 33'b0101100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2451] = 33'b0100000101100000_0_0_xx_110_001_xxx_1_x_xx;
      patterns[2452] = 33'b0100100101100000_1_0_xx_110_001_xxx_1_x_xx;
      patterns[2453] = 33'b0100100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2454] = 33'b0000000111000101_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2455] = 33'b0000100111000101_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2456] = 33'b0000100111000101_0_0_00_000_000_000_0_0_00;
      patterns[2457] = 33'b1000000101100101_0_1_00_110_101_001_0_x_00;
      patterns[2458] = 33'b1000100101100101_1_1_00_110_101_001_0_x_00;
      patterns[2459] = 33'b1000100101100101_0_0_00_000_000_000_0_0_00;
      patterns[2460] = 33'b1001000101100101_0_1_01_110_101_001_0_x_00;
      patterns[2461] = 33'b1001100101100101_1_1_01_110_101_001_0_x_00;
      patterns[2462] = 33'b1001100101100101_0_0_00_000_000_000_0_0_00;
      patterns[2463] = 33'b1010000101100101_0_1_10_110_101_001_0_x_00;
      patterns[2464] = 33'b1010100101100101_1_1_10_110_101_001_0_x_00;
      patterns[2465] = 33'b1010100101100101_0_0_00_000_000_000_0_0_00;
      patterns[2466] = 33'b1011000101100101_0_1_11_110_101_001_0_x_00;
      patterns[2467] = 33'b1011100101100101_1_1_11_110_101_001_0_x_00;
      patterns[2468] = 33'b1011100101100101_0_0_00_000_000_000_0_0_00;
      patterns[2469] = 33'b0101000101100000_0_1_xx_110_xxx_001_0_1_01;
      patterns[2470] = 33'b0101100101100000_1_1_xx_110_xxx_001_0_1_01;
      patterns[2471] = 33'b0101100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2472] = 33'b0100000101100000_0_0_xx_110_001_xxx_1_x_xx;
      patterns[2473] = 33'b0100100101100000_1_0_xx_110_001_xxx_1_x_xx;
      patterns[2474] = 33'b0100100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2475] = 33'b0000000110111011_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2476] = 33'b0000100110111011_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2477] = 33'b0000100110111011_0_0_00_000_000_000_0_0_00;
      patterns[2478] = 33'b1000000101100110_0_1_00_110_110_001_0_x_00;
      patterns[2479] = 33'b1000100101100110_1_1_00_110_110_001_0_x_00;
      patterns[2480] = 33'b1000100101100110_0_0_00_000_000_000_0_0_00;
      patterns[2481] = 33'b1001000101100110_0_1_01_110_110_001_0_x_00;
      patterns[2482] = 33'b1001100101100110_1_1_01_110_110_001_0_x_00;
      patterns[2483] = 33'b1001100101100110_0_0_00_000_000_000_0_0_00;
      patterns[2484] = 33'b1010000101100110_0_1_10_110_110_001_0_x_00;
      patterns[2485] = 33'b1010100101100110_1_1_10_110_110_001_0_x_00;
      patterns[2486] = 33'b1010100101100110_0_0_00_000_000_000_0_0_00;
      patterns[2487] = 33'b1011000101100110_0_1_11_110_110_001_0_x_00;
      patterns[2488] = 33'b1011100101100110_1_1_11_110_110_001_0_x_00;
      patterns[2489] = 33'b1011100101100110_0_0_00_000_000_000_0_0_00;
      patterns[2490] = 33'b0101000101100000_0_1_xx_110_xxx_001_0_1_01;
      patterns[2491] = 33'b0101100101100000_1_1_xx_110_xxx_001_0_1_01;
      patterns[2492] = 33'b0101100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2493] = 33'b0100000101100000_0_0_xx_110_001_xxx_1_x_xx;
      patterns[2494] = 33'b0100100101100000_1_0_xx_110_001_xxx_1_x_xx;
      patterns[2495] = 33'b0100100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2496] = 33'b0000000100101110_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2497] = 33'b0000100100101110_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2498] = 33'b0000100100101110_0_0_00_000_000_000_0_0_00;
      patterns[2499] = 33'b1000000101100111_0_1_00_110_111_001_0_x_00;
      patterns[2500] = 33'b1000100101100111_1_1_00_110_111_001_0_x_00;
      patterns[2501] = 33'b1000100101100111_0_0_00_000_000_000_0_0_00;
      patterns[2502] = 33'b1001000101100111_0_1_01_110_111_001_0_x_00;
      patterns[2503] = 33'b1001100101100111_1_1_01_110_111_001_0_x_00;
      patterns[2504] = 33'b1001100101100111_0_0_00_000_000_000_0_0_00;
      patterns[2505] = 33'b1010000101100111_0_1_10_110_111_001_0_x_00;
      patterns[2506] = 33'b1010100101100111_1_1_10_110_111_001_0_x_00;
      patterns[2507] = 33'b1010100101100111_0_0_00_000_000_000_0_0_00;
      patterns[2508] = 33'b1011000101100111_0_1_11_110_111_001_0_x_00;
      patterns[2509] = 33'b1011100101100111_1_1_11_110_111_001_0_x_00;
      patterns[2510] = 33'b1011100101100111_0_0_00_000_000_000_0_0_00;
      patterns[2511] = 33'b0101000101100000_0_1_xx_110_xxx_001_0_1_01;
      patterns[2512] = 33'b0101100101100000_1_1_xx_110_xxx_001_0_1_01;
      patterns[2513] = 33'b0101100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2514] = 33'b0100000101100000_0_0_xx_110_001_xxx_1_x_xx;
      patterns[2515] = 33'b0100100101100000_1_0_xx_110_001_xxx_1_x_xx;
      patterns[2516] = 33'b0100100101100000_0_0_00_000_000_000_0_0_00;
      patterns[2517] = 33'b0000000100000000_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2518] = 33'b0000100100000000_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2519] = 33'b0000100100000000_0_0_00_000_000_000_0_0_00;
      patterns[2520] = 33'b1000000101110000_0_1_00_111_000_001_0_x_00;
      patterns[2521] = 33'b1000100101110000_1_1_00_111_000_001_0_x_00;
      patterns[2522] = 33'b1000100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2523] = 33'b1001000101110000_0_1_01_111_000_001_0_x_00;
      patterns[2524] = 33'b1001100101110000_1_1_01_111_000_001_0_x_00;
      patterns[2525] = 33'b1001100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2526] = 33'b1010000101110000_0_1_10_111_000_001_0_x_00;
      patterns[2527] = 33'b1010100101110000_1_1_10_111_000_001_0_x_00;
      patterns[2528] = 33'b1010100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2529] = 33'b1011000101110000_0_1_11_111_000_001_0_x_00;
      patterns[2530] = 33'b1011100101110000_1_1_11_111_000_001_0_x_00;
      patterns[2531] = 33'b1011100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2532] = 33'b0101000101110000_0_1_xx_111_xxx_001_0_1_01;
      patterns[2533] = 33'b0101100101110000_1_1_xx_111_xxx_001_0_1_01;
      patterns[2534] = 33'b0101100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2535] = 33'b0100000101110000_0_0_xx_111_001_xxx_1_x_xx;
      patterns[2536] = 33'b0100100101110000_1_0_xx_111_001_xxx_1_x_xx;
      patterns[2537] = 33'b0100100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2538] = 33'b0000000100000110_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2539] = 33'b0000100100000110_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2540] = 33'b0000100100000110_0_0_00_000_000_000_0_0_00;
      patterns[2541] = 33'b1000000101110001_0_1_00_111_001_001_0_x_00;
      patterns[2542] = 33'b1000100101110001_1_1_00_111_001_001_0_x_00;
      patterns[2543] = 33'b1000100101110001_0_0_00_000_000_000_0_0_00;
      patterns[2544] = 33'b1001000101110001_0_1_01_111_001_001_0_x_00;
      patterns[2545] = 33'b1001100101110001_1_1_01_111_001_001_0_x_00;
      patterns[2546] = 33'b1001100101110001_0_0_00_000_000_000_0_0_00;
      patterns[2547] = 33'b1010000101110001_0_1_10_111_001_001_0_x_00;
      patterns[2548] = 33'b1010100101110001_1_1_10_111_001_001_0_x_00;
      patterns[2549] = 33'b1010100101110001_0_0_00_000_000_000_0_0_00;
      patterns[2550] = 33'b1011000101110001_0_1_11_111_001_001_0_x_00;
      patterns[2551] = 33'b1011100101110001_1_1_11_111_001_001_0_x_00;
      patterns[2552] = 33'b1011100101110001_0_0_00_000_000_000_0_0_00;
      patterns[2553] = 33'b0101000101110000_0_1_xx_111_xxx_001_0_1_01;
      patterns[2554] = 33'b0101100101110000_1_1_xx_111_xxx_001_0_1_01;
      patterns[2555] = 33'b0101100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2556] = 33'b0100000101110000_0_0_xx_111_001_xxx_1_x_xx;
      patterns[2557] = 33'b0100100101110000_1_0_xx_111_001_xxx_1_x_xx;
      patterns[2558] = 33'b0100100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2559] = 33'b0000000110000110_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2560] = 33'b0000100110000110_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2561] = 33'b0000100110000110_0_0_00_000_000_000_0_0_00;
      patterns[2562] = 33'b1000000101110010_0_1_00_111_010_001_0_x_00;
      patterns[2563] = 33'b1000100101110010_1_1_00_111_010_001_0_x_00;
      patterns[2564] = 33'b1000100101110010_0_0_00_000_000_000_0_0_00;
      patterns[2565] = 33'b1001000101110010_0_1_01_111_010_001_0_x_00;
      patterns[2566] = 33'b1001100101110010_1_1_01_111_010_001_0_x_00;
      patterns[2567] = 33'b1001100101110010_0_0_00_000_000_000_0_0_00;
      patterns[2568] = 33'b1010000101110010_0_1_10_111_010_001_0_x_00;
      patterns[2569] = 33'b1010100101110010_1_1_10_111_010_001_0_x_00;
      patterns[2570] = 33'b1010100101110010_0_0_00_000_000_000_0_0_00;
      patterns[2571] = 33'b1011000101110010_0_1_11_111_010_001_0_x_00;
      patterns[2572] = 33'b1011100101110010_1_1_11_111_010_001_0_x_00;
      patterns[2573] = 33'b1011100101110010_0_0_00_000_000_000_0_0_00;
      patterns[2574] = 33'b0101000101110000_0_1_xx_111_xxx_001_0_1_01;
      patterns[2575] = 33'b0101100101110000_1_1_xx_111_xxx_001_0_1_01;
      patterns[2576] = 33'b0101100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2577] = 33'b0100000101110000_0_0_xx_111_001_xxx_1_x_xx;
      patterns[2578] = 33'b0100100101110000_1_0_xx_111_001_xxx_1_x_xx;
      patterns[2579] = 33'b0100100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2580] = 33'b0000000111111110_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2581] = 33'b0000100111111110_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2582] = 33'b0000100111111110_0_0_00_000_000_000_0_0_00;
      patterns[2583] = 33'b1000000101110011_0_1_00_111_011_001_0_x_00;
      patterns[2584] = 33'b1000100101110011_1_1_00_111_011_001_0_x_00;
      patterns[2585] = 33'b1000100101110011_0_0_00_000_000_000_0_0_00;
      patterns[2586] = 33'b1001000101110011_0_1_01_111_011_001_0_x_00;
      patterns[2587] = 33'b1001100101110011_1_1_01_111_011_001_0_x_00;
      patterns[2588] = 33'b1001100101110011_0_0_00_000_000_000_0_0_00;
      patterns[2589] = 33'b1010000101110011_0_1_10_111_011_001_0_x_00;
      patterns[2590] = 33'b1010100101110011_1_1_10_111_011_001_0_x_00;
      patterns[2591] = 33'b1010100101110011_0_0_00_000_000_000_0_0_00;
      patterns[2592] = 33'b1011000101110011_0_1_11_111_011_001_0_x_00;
      patterns[2593] = 33'b1011100101110011_1_1_11_111_011_001_0_x_00;
      patterns[2594] = 33'b1011100101110011_0_0_00_000_000_000_0_0_00;
      patterns[2595] = 33'b0101000101110000_0_1_xx_111_xxx_001_0_1_01;
      patterns[2596] = 33'b0101100101110000_1_1_xx_111_xxx_001_0_1_01;
      patterns[2597] = 33'b0101100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2598] = 33'b0100000101110000_0_0_xx_111_001_xxx_1_x_xx;
      patterns[2599] = 33'b0100100101110000_1_0_xx_111_001_xxx_1_x_xx;
      patterns[2600] = 33'b0100100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2601] = 33'b0000000110011010_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2602] = 33'b0000100110011010_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2603] = 33'b0000100110011010_0_0_00_000_000_000_0_0_00;
      patterns[2604] = 33'b1000000101110100_0_1_00_111_100_001_0_x_00;
      patterns[2605] = 33'b1000100101110100_1_1_00_111_100_001_0_x_00;
      patterns[2606] = 33'b1000100101110100_0_0_00_000_000_000_0_0_00;
      patterns[2607] = 33'b1001000101110100_0_1_01_111_100_001_0_x_00;
      patterns[2608] = 33'b1001100101110100_1_1_01_111_100_001_0_x_00;
      patterns[2609] = 33'b1001100101110100_0_0_00_000_000_000_0_0_00;
      patterns[2610] = 33'b1010000101110100_0_1_10_111_100_001_0_x_00;
      patterns[2611] = 33'b1010100101110100_1_1_10_111_100_001_0_x_00;
      patterns[2612] = 33'b1010100101110100_0_0_00_000_000_000_0_0_00;
      patterns[2613] = 33'b1011000101110100_0_1_11_111_100_001_0_x_00;
      patterns[2614] = 33'b1011100101110100_1_1_11_111_100_001_0_x_00;
      patterns[2615] = 33'b1011100101110100_0_0_00_000_000_000_0_0_00;
      patterns[2616] = 33'b0101000101110000_0_1_xx_111_xxx_001_0_1_01;
      patterns[2617] = 33'b0101100101110000_1_1_xx_111_xxx_001_0_1_01;
      patterns[2618] = 33'b0101100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2619] = 33'b0100000101110000_0_0_xx_111_001_xxx_1_x_xx;
      patterns[2620] = 33'b0100100101110000_1_0_xx_111_001_xxx_1_x_xx;
      patterns[2621] = 33'b0100100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2622] = 33'b0000000100000100_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2623] = 33'b0000100100000100_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2624] = 33'b0000100100000100_0_0_00_000_000_000_0_0_00;
      patterns[2625] = 33'b1000000101110101_0_1_00_111_101_001_0_x_00;
      patterns[2626] = 33'b1000100101110101_1_1_00_111_101_001_0_x_00;
      patterns[2627] = 33'b1000100101110101_0_0_00_000_000_000_0_0_00;
      patterns[2628] = 33'b1001000101110101_0_1_01_111_101_001_0_x_00;
      patterns[2629] = 33'b1001100101110101_1_1_01_111_101_001_0_x_00;
      patterns[2630] = 33'b1001100101110101_0_0_00_000_000_000_0_0_00;
      patterns[2631] = 33'b1010000101110101_0_1_10_111_101_001_0_x_00;
      patterns[2632] = 33'b1010100101110101_1_1_10_111_101_001_0_x_00;
      patterns[2633] = 33'b1010100101110101_0_0_00_000_000_000_0_0_00;
      patterns[2634] = 33'b1011000101110101_0_1_11_111_101_001_0_x_00;
      patterns[2635] = 33'b1011100101110101_1_1_11_111_101_001_0_x_00;
      patterns[2636] = 33'b1011100101110101_0_0_00_000_000_000_0_0_00;
      patterns[2637] = 33'b0101000101110000_0_1_xx_111_xxx_001_0_1_01;
      patterns[2638] = 33'b0101100101110000_1_1_xx_111_xxx_001_0_1_01;
      patterns[2639] = 33'b0101100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2640] = 33'b0100000101110000_0_0_xx_111_001_xxx_1_x_xx;
      patterns[2641] = 33'b0100100101110000_1_0_xx_111_001_xxx_1_x_xx;
      patterns[2642] = 33'b0100100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2643] = 33'b0000000100110001_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2644] = 33'b0000100100110001_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2645] = 33'b0000100100110001_0_0_00_000_000_000_0_0_00;
      patterns[2646] = 33'b1000000101110110_0_1_00_111_110_001_0_x_00;
      patterns[2647] = 33'b1000100101110110_1_1_00_111_110_001_0_x_00;
      patterns[2648] = 33'b1000100101110110_0_0_00_000_000_000_0_0_00;
      patterns[2649] = 33'b1001000101110110_0_1_01_111_110_001_0_x_00;
      patterns[2650] = 33'b1001100101110110_1_1_01_111_110_001_0_x_00;
      patterns[2651] = 33'b1001100101110110_0_0_00_000_000_000_0_0_00;
      patterns[2652] = 33'b1010000101110110_0_1_10_111_110_001_0_x_00;
      patterns[2653] = 33'b1010100101110110_1_1_10_111_110_001_0_x_00;
      patterns[2654] = 33'b1010100101110110_0_0_00_000_000_000_0_0_00;
      patterns[2655] = 33'b1011000101110110_0_1_11_111_110_001_0_x_00;
      patterns[2656] = 33'b1011100101110110_1_1_11_111_110_001_0_x_00;
      patterns[2657] = 33'b1011100101110110_0_0_00_000_000_000_0_0_00;
      patterns[2658] = 33'b0101000101110000_0_1_xx_111_xxx_001_0_1_01;
      patterns[2659] = 33'b0101100101110000_1_1_xx_111_xxx_001_0_1_01;
      patterns[2660] = 33'b0101100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2661] = 33'b0100000101110000_0_0_xx_111_001_xxx_1_x_xx;
      patterns[2662] = 33'b0100100101110000_1_0_xx_111_001_xxx_1_x_xx;
      patterns[2663] = 33'b0100100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2664] = 33'b0000000110011100_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2665] = 33'b0000100110011100_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2666] = 33'b0000100110011100_0_0_00_000_000_000_0_0_00;
      patterns[2667] = 33'b1000000101110111_0_1_00_111_111_001_0_x_00;
      patterns[2668] = 33'b1000100101110111_1_1_00_111_111_001_0_x_00;
      patterns[2669] = 33'b1000100101110111_0_0_00_000_000_000_0_0_00;
      patterns[2670] = 33'b1001000101110111_0_1_01_111_111_001_0_x_00;
      patterns[2671] = 33'b1001100101110111_1_1_01_111_111_001_0_x_00;
      patterns[2672] = 33'b1001100101110111_0_0_00_000_000_000_0_0_00;
      patterns[2673] = 33'b1010000101110111_0_1_10_111_111_001_0_x_00;
      patterns[2674] = 33'b1010100101110111_1_1_10_111_111_001_0_x_00;
      patterns[2675] = 33'b1010100101110111_0_0_00_000_000_000_0_0_00;
      patterns[2676] = 33'b1011000101110111_0_1_11_111_111_001_0_x_00;
      patterns[2677] = 33'b1011100101110111_1_1_11_111_111_001_0_x_00;
      patterns[2678] = 33'b1011100101110111_0_0_00_000_000_000_0_0_00;
      patterns[2679] = 33'b0101000101110000_0_1_xx_111_xxx_001_0_1_01;
      patterns[2680] = 33'b0101100101110000_1_1_xx_111_xxx_001_0_1_01;
      patterns[2681] = 33'b0101100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2682] = 33'b0100000101110000_0_0_xx_111_001_xxx_1_x_xx;
      patterns[2683] = 33'b0100100101110000_1_0_xx_111_001_xxx_1_x_xx;
      patterns[2684] = 33'b0100100101110000_0_0_00_000_000_000_0_0_00;
      patterns[2685] = 33'b0000000101111110_0_1_xx_xxx_xxx_001_0_x_10;
      patterns[2686] = 33'b0000100101111110_1_1_xx_xxx_xxx_001_0_x_10;
      patterns[2687] = 33'b0000100101111110_0_0_00_000_000_000_0_0_00;
      patterns[2688] = 33'b1000001000000000_0_1_00_000_000_010_0_x_00;
      patterns[2689] = 33'b1000101000000000_1_1_00_000_000_010_0_x_00;
      patterns[2690] = 33'b1000101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2691] = 33'b1001001000000000_0_1_01_000_000_010_0_x_00;
      patterns[2692] = 33'b1001101000000000_1_1_01_000_000_010_0_x_00;
      patterns[2693] = 33'b1001101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2694] = 33'b1010001000000000_0_1_10_000_000_010_0_x_00;
      patterns[2695] = 33'b1010101000000000_1_1_10_000_000_010_0_x_00;
      patterns[2696] = 33'b1010101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2697] = 33'b1011001000000000_0_1_11_000_000_010_0_x_00;
      patterns[2698] = 33'b1011101000000000_1_1_11_000_000_010_0_x_00;
      patterns[2699] = 33'b1011101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2700] = 33'b0101001000000000_0_1_xx_000_xxx_010_0_1_01;
      patterns[2701] = 33'b0101101000000000_1_1_xx_000_xxx_010_0_1_01;
      patterns[2702] = 33'b0101101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2703] = 33'b0100001000000000_0_0_xx_000_010_xxx_1_x_xx;
      patterns[2704] = 33'b0100101000000000_1_0_xx_000_010_xxx_1_x_xx;
      patterns[2705] = 33'b0100101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2706] = 33'b0000001001110100_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[2707] = 33'b0000101001110100_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[2708] = 33'b0000101001110100_0_0_00_000_000_000_0_0_00;
      patterns[2709] = 33'b1000001000000001_0_1_00_000_001_010_0_x_00;
      patterns[2710] = 33'b1000101000000001_1_1_00_000_001_010_0_x_00;
      patterns[2711] = 33'b1000101000000001_0_0_00_000_000_000_0_0_00;
      patterns[2712] = 33'b1001001000000001_0_1_01_000_001_010_0_x_00;
      patterns[2713] = 33'b1001101000000001_1_1_01_000_001_010_0_x_00;
      patterns[2714] = 33'b1001101000000001_0_0_00_000_000_000_0_0_00;
      patterns[2715] = 33'b1010001000000001_0_1_10_000_001_010_0_x_00;
      patterns[2716] = 33'b1010101000000001_1_1_10_000_001_010_0_x_00;
      patterns[2717] = 33'b1010101000000001_0_0_00_000_000_000_0_0_00;
      patterns[2718] = 33'b1011001000000001_0_1_11_000_001_010_0_x_00;
      patterns[2719] = 33'b1011101000000001_1_1_11_000_001_010_0_x_00;
      patterns[2720] = 33'b1011101000000001_0_0_00_000_000_000_0_0_00;
      patterns[2721] = 33'b0101001000000000_0_1_xx_000_xxx_010_0_1_01;
      patterns[2722] = 33'b0101101000000000_1_1_xx_000_xxx_010_0_1_01;
      patterns[2723] = 33'b0101101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2724] = 33'b0100001000000000_0_0_xx_000_010_xxx_1_x_xx;
      patterns[2725] = 33'b0100101000000000_1_0_xx_000_010_xxx_1_x_xx;
      patterns[2726] = 33'b0100101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2727] = 33'b0000001001110001_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[2728] = 33'b0000101001110001_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[2729] = 33'b0000101001110001_0_0_00_000_000_000_0_0_00;
      patterns[2730] = 33'b1000001000000010_0_1_00_000_010_010_0_x_00;
      patterns[2731] = 33'b1000101000000010_1_1_00_000_010_010_0_x_00;
      patterns[2732] = 33'b1000101000000010_0_0_00_000_000_000_0_0_00;
      patterns[2733] = 33'b1001001000000010_0_1_01_000_010_010_0_x_00;
      patterns[2734] = 33'b1001101000000010_1_1_01_000_010_010_0_x_00;
      patterns[2735] = 33'b1001101000000010_0_0_00_000_000_000_0_0_00;
      patterns[2736] = 33'b1010001000000010_0_1_10_000_010_010_0_x_00;
      patterns[2737] = 33'b1010101000000010_1_1_10_000_010_010_0_x_00;
      patterns[2738] = 33'b1010101000000010_0_0_00_000_000_000_0_0_00;
      patterns[2739] = 33'b1011001000000010_0_1_11_000_010_010_0_x_00;
      patterns[2740] = 33'b1011101000000010_1_1_11_000_010_010_0_x_00;
      patterns[2741] = 33'b1011101000000010_0_0_00_000_000_000_0_0_00;
      patterns[2742] = 33'b0101001000000000_0_1_xx_000_xxx_010_0_1_01;
      patterns[2743] = 33'b0101101000000000_1_1_xx_000_xxx_010_0_1_01;
      patterns[2744] = 33'b0101101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2745] = 33'b0100001000000000_0_0_xx_000_010_xxx_1_x_xx;
      patterns[2746] = 33'b0100101000000000_1_0_xx_000_010_xxx_1_x_xx;
      patterns[2747] = 33'b0100101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2748] = 33'b0000001010110000_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[2749] = 33'b0000101010110000_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[2750] = 33'b0000101010110000_0_0_00_000_000_000_0_0_00;
      patterns[2751] = 33'b1000001000000011_0_1_00_000_011_010_0_x_00;
      patterns[2752] = 33'b1000101000000011_1_1_00_000_011_010_0_x_00;
      patterns[2753] = 33'b1000101000000011_0_0_00_000_000_000_0_0_00;
      patterns[2754] = 33'b1001001000000011_0_1_01_000_011_010_0_x_00;
      patterns[2755] = 33'b1001101000000011_1_1_01_000_011_010_0_x_00;
      patterns[2756] = 33'b1001101000000011_0_0_00_000_000_000_0_0_00;
      patterns[2757] = 33'b1010001000000011_0_1_10_000_011_010_0_x_00;
      patterns[2758] = 33'b1010101000000011_1_1_10_000_011_010_0_x_00;
      patterns[2759] = 33'b1010101000000011_0_0_00_000_000_000_0_0_00;
      patterns[2760] = 33'b1011001000000011_0_1_11_000_011_010_0_x_00;
      patterns[2761] = 33'b1011101000000011_1_1_11_000_011_010_0_x_00;
      patterns[2762] = 33'b1011101000000011_0_0_00_000_000_000_0_0_00;
      patterns[2763] = 33'b0101001000000000_0_1_xx_000_xxx_010_0_1_01;
      patterns[2764] = 33'b0101101000000000_1_1_xx_000_xxx_010_0_1_01;
      patterns[2765] = 33'b0101101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2766] = 33'b0100001000000000_0_0_xx_000_010_xxx_1_x_xx;
      patterns[2767] = 33'b0100101000000000_1_0_xx_000_010_xxx_1_x_xx;
      patterns[2768] = 33'b0100101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2769] = 33'b0000001010000000_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[2770] = 33'b0000101010000000_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[2771] = 33'b0000101010000000_0_0_00_000_000_000_0_0_00;
      patterns[2772] = 33'b1000001000000100_0_1_00_000_100_010_0_x_00;
      patterns[2773] = 33'b1000101000000100_1_1_00_000_100_010_0_x_00;
      patterns[2774] = 33'b1000101000000100_0_0_00_000_000_000_0_0_00;
      patterns[2775] = 33'b1001001000000100_0_1_01_000_100_010_0_x_00;
      patterns[2776] = 33'b1001101000000100_1_1_01_000_100_010_0_x_00;
      patterns[2777] = 33'b1001101000000100_0_0_00_000_000_000_0_0_00;
      patterns[2778] = 33'b1010001000000100_0_1_10_000_100_010_0_x_00;
      patterns[2779] = 33'b1010101000000100_1_1_10_000_100_010_0_x_00;
      patterns[2780] = 33'b1010101000000100_0_0_00_000_000_000_0_0_00;
      patterns[2781] = 33'b1011001000000100_0_1_11_000_100_010_0_x_00;
      patterns[2782] = 33'b1011101000000100_1_1_11_000_100_010_0_x_00;
      patterns[2783] = 33'b1011101000000100_0_0_00_000_000_000_0_0_00;
      patterns[2784] = 33'b0101001000000000_0_1_xx_000_xxx_010_0_1_01;
      patterns[2785] = 33'b0101101000000000_1_1_xx_000_xxx_010_0_1_01;
      patterns[2786] = 33'b0101101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2787] = 33'b0100001000000000_0_0_xx_000_010_xxx_1_x_xx;
      patterns[2788] = 33'b0100101000000000_1_0_xx_000_010_xxx_1_x_xx;
      patterns[2789] = 33'b0100101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2790] = 33'b0000001000000110_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[2791] = 33'b0000101000000110_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[2792] = 33'b0000101000000110_0_0_00_000_000_000_0_0_00;
      patterns[2793] = 33'b1000001000000101_0_1_00_000_101_010_0_x_00;
      patterns[2794] = 33'b1000101000000101_1_1_00_000_101_010_0_x_00;
      patterns[2795] = 33'b1000101000000101_0_0_00_000_000_000_0_0_00;
      patterns[2796] = 33'b1001001000000101_0_1_01_000_101_010_0_x_00;
      patterns[2797] = 33'b1001101000000101_1_1_01_000_101_010_0_x_00;
      patterns[2798] = 33'b1001101000000101_0_0_00_000_000_000_0_0_00;
      patterns[2799] = 33'b1010001000000101_0_1_10_000_101_010_0_x_00;
      patterns[2800] = 33'b1010101000000101_1_1_10_000_101_010_0_x_00;
      patterns[2801] = 33'b1010101000000101_0_0_00_000_000_000_0_0_00;
      patterns[2802] = 33'b1011001000000101_0_1_11_000_101_010_0_x_00;
      patterns[2803] = 33'b1011101000000101_1_1_11_000_101_010_0_x_00;
      patterns[2804] = 33'b1011101000000101_0_0_00_000_000_000_0_0_00;
      patterns[2805] = 33'b0101001000000000_0_1_xx_000_xxx_010_0_1_01;
      patterns[2806] = 33'b0101101000000000_1_1_xx_000_xxx_010_0_1_01;
      patterns[2807] = 33'b0101101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2808] = 33'b0100001000000000_0_0_xx_000_010_xxx_1_x_xx;
      patterns[2809] = 33'b0100101000000000_1_0_xx_000_010_xxx_1_x_xx;
      patterns[2810] = 33'b0100101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2811] = 33'b0000001000001111_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[2812] = 33'b0000101000001111_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[2813] = 33'b0000101000001111_0_0_00_000_000_000_0_0_00;
      patterns[2814] = 33'b1000001000000110_0_1_00_000_110_010_0_x_00;
      patterns[2815] = 33'b1000101000000110_1_1_00_000_110_010_0_x_00;
      patterns[2816] = 33'b1000101000000110_0_0_00_000_000_000_0_0_00;
      patterns[2817] = 33'b1001001000000110_0_1_01_000_110_010_0_x_00;
      patterns[2818] = 33'b1001101000000110_1_1_01_000_110_010_0_x_00;
      patterns[2819] = 33'b1001101000000110_0_0_00_000_000_000_0_0_00;
      patterns[2820] = 33'b1010001000000110_0_1_10_000_110_010_0_x_00;
      patterns[2821] = 33'b1010101000000110_1_1_10_000_110_010_0_x_00;
      patterns[2822] = 33'b1010101000000110_0_0_00_000_000_000_0_0_00;
      patterns[2823] = 33'b1011001000000110_0_1_11_000_110_010_0_x_00;
      patterns[2824] = 33'b1011101000000110_1_1_11_000_110_010_0_x_00;
      patterns[2825] = 33'b1011101000000110_0_0_00_000_000_000_0_0_00;
      patterns[2826] = 33'b0101001000000000_0_1_xx_000_xxx_010_0_1_01;
      patterns[2827] = 33'b0101101000000000_1_1_xx_000_xxx_010_0_1_01;
      patterns[2828] = 33'b0101101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2829] = 33'b0100001000000000_0_0_xx_000_010_xxx_1_x_xx;
      patterns[2830] = 33'b0100101000000000_1_0_xx_000_010_xxx_1_x_xx;
      patterns[2831] = 33'b0100101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2832] = 33'b0000001010100011_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[2833] = 33'b0000101010100011_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[2834] = 33'b0000101010100011_0_0_00_000_000_000_0_0_00;
      patterns[2835] = 33'b1000001000000111_0_1_00_000_111_010_0_x_00;
      patterns[2836] = 33'b1000101000000111_1_1_00_000_111_010_0_x_00;
      patterns[2837] = 33'b1000101000000111_0_0_00_000_000_000_0_0_00;
      patterns[2838] = 33'b1001001000000111_0_1_01_000_111_010_0_x_00;
      patterns[2839] = 33'b1001101000000111_1_1_01_000_111_010_0_x_00;
      patterns[2840] = 33'b1001101000000111_0_0_00_000_000_000_0_0_00;
      patterns[2841] = 33'b1010001000000111_0_1_10_000_111_010_0_x_00;
      patterns[2842] = 33'b1010101000000111_1_1_10_000_111_010_0_x_00;
      patterns[2843] = 33'b1010101000000111_0_0_00_000_000_000_0_0_00;
      patterns[2844] = 33'b1011001000000111_0_1_11_000_111_010_0_x_00;
      patterns[2845] = 33'b1011101000000111_1_1_11_000_111_010_0_x_00;
      patterns[2846] = 33'b1011101000000111_0_0_00_000_000_000_0_0_00;
      patterns[2847] = 33'b0101001000000000_0_1_xx_000_xxx_010_0_1_01;
      patterns[2848] = 33'b0101101000000000_1_1_xx_000_xxx_010_0_1_01;
      patterns[2849] = 33'b0101101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2850] = 33'b0100001000000000_0_0_xx_000_010_xxx_1_x_xx;
      patterns[2851] = 33'b0100101000000000_1_0_xx_000_010_xxx_1_x_xx;
      patterns[2852] = 33'b0100101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2853] = 33'b0000001000001101_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[2854] = 33'b0000101000001101_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[2855] = 33'b0000101000001101_0_0_00_000_000_000_0_0_00;
      patterns[2856] = 33'b1000001000010000_0_1_00_001_000_010_0_x_00;
      patterns[2857] = 33'b1000101000010000_1_1_00_001_000_010_0_x_00;
      patterns[2858] = 33'b1000101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2859] = 33'b1001001000010000_0_1_01_001_000_010_0_x_00;
      patterns[2860] = 33'b1001101000010000_1_1_01_001_000_010_0_x_00;
      patterns[2861] = 33'b1001101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2862] = 33'b1010001000010000_0_1_10_001_000_010_0_x_00;
      patterns[2863] = 33'b1010101000010000_1_1_10_001_000_010_0_x_00;
      patterns[2864] = 33'b1010101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2865] = 33'b1011001000010000_0_1_11_001_000_010_0_x_00;
      patterns[2866] = 33'b1011101000010000_1_1_11_001_000_010_0_x_00;
      patterns[2867] = 33'b1011101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2868] = 33'b0101001000010000_0_1_xx_001_xxx_010_0_1_01;
      patterns[2869] = 33'b0101101000010000_1_1_xx_001_xxx_010_0_1_01;
      patterns[2870] = 33'b0101101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2871] = 33'b0100001000010000_0_0_xx_001_010_xxx_1_x_xx;
      patterns[2872] = 33'b0100101000010000_1_0_xx_001_010_xxx_1_x_xx;
      patterns[2873] = 33'b0100101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2874] = 33'b0000001011001110_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[2875] = 33'b0000101011001110_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[2876] = 33'b0000101011001110_0_0_00_000_000_000_0_0_00;
      patterns[2877] = 33'b1000001000010001_0_1_00_001_001_010_0_x_00;
      patterns[2878] = 33'b1000101000010001_1_1_00_001_001_010_0_x_00;
      patterns[2879] = 33'b1000101000010001_0_0_00_000_000_000_0_0_00;
      patterns[2880] = 33'b1001001000010001_0_1_01_001_001_010_0_x_00;
      patterns[2881] = 33'b1001101000010001_1_1_01_001_001_010_0_x_00;
      patterns[2882] = 33'b1001101000010001_0_0_00_000_000_000_0_0_00;
      patterns[2883] = 33'b1010001000010001_0_1_10_001_001_010_0_x_00;
      patterns[2884] = 33'b1010101000010001_1_1_10_001_001_010_0_x_00;
      patterns[2885] = 33'b1010101000010001_0_0_00_000_000_000_0_0_00;
      patterns[2886] = 33'b1011001000010001_0_1_11_001_001_010_0_x_00;
      patterns[2887] = 33'b1011101000010001_1_1_11_001_001_010_0_x_00;
      patterns[2888] = 33'b1011101000010001_0_0_00_000_000_000_0_0_00;
      patterns[2889] = 33'b0101001000010000_0_1_xx_001_xxx_010_0_1_01;
      patterns[2890] = 33'b0101101000010000_1_1_xx_001_xxx_010_0_1_01;
      patterns[2891] = 33'b0101101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2892] = 33'b0100001000010000_0_0_xx_001_010_xxx_1_x_xx;
      patterns[2893] = 33'b0100101000010000_1_0_xx_001_010_xxx_1_x_xx;
      patterns[2894] = 33'b0100101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2895] = 33'b0000001010101100_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[2896] = 33'b0000101010101100_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[2897] = 33'b0000101010101100_0_0_00_000_000_000_0_0_00;
      patterns[2898] = 33'b1000001000010010_0_1_00_001_010_010_0_x_00;
      patterns[2899] = 33'b1000101000010010_1_1_00_001_010_010_0_x_00;
      patterns[2900] = 33'b1000101000010010_0_0_00_000_000_000_0_0_00;
      patterns[2901] = 33'b1001001000010010_0_1_01_001_010_010_0_x_00;
      patterns[2902] = 33'b1001101000010010_1_1_01_001_010_010_0_x_00;
      patterns[2903] = 33'b1001101000010010_0_0_00_000_000_000_0_0_00;
      patterns[2904] = 33'b1010001000010010_0_1_10_001_010_010_0_x_00;
      patterns[2905] = 33'b1010101000010010_1_1_10_001_010_010_0_x_00;
      patterns[2906] = 33'b1010101000010010_0_0_00_000_000_000_0_0_00;
      patterns[2907] = 33'b1011001000010010_0_1_11_001_010_010_0_x_00;
      patterns[2908] = 33'b1011101000010010_1_1_11_001_010_010_0_x_00;
      patterns[2909] = 33'b1011101000010010_0_0_00_000_000_000_0_0_00;
      patterns[2910] = 33'b0101001000010000_0_1_xx_001_xxx_010_0_1_01;
      patterns[2911] = 33'b0101101000010000_1_1_xx_001_xxx_010_0_1_01;
      patterns[2912] = 33'b0101101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2913] = 33'b0100001000010000_0_0_xx_001_010_xxx_1_x_xx;
      patterns[2914] = 33'b0100101000010000_1_0_xx_001_010_xxx_1_x_xx;
      patterns[2915] = 33'b0100101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2916] = 33'b0000001011100101_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[2917] = 33'b0000101011100101_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[2918] = 33'b0000101011100101_0_0_00_000_000_000_0_0_00;
      patterns[2919] = 33'b1000001000010011_0_1_00_001_011_010_0_x_00;
      patterns[2920] = 33'b1000101000010011_1_1_00_001_011_010_0_x_00;
      patterns[2921] = 33'b1000101000010011_0_0_00_000_000_000_0_0_00;
      patterns[2922] = 33'b1001001000010011_0_1_01_001_011_010_0_x_00;
      patterns[2923] = 33'b1001101000010011_1_1_01_001_011_010_0_x_00;
      patterns[2924] = 33'b1001101000010011_0_0_00_000_000_000_0_0_00;
      patterns[2925] = 33'b1010001000010011_0_1_10_001_011_010_0_x_00;
      patterns[2926] = 33'b1010101000010011_1_1_10_001_011_010_0_x_00;
      patterns[2927] = 33'b1010101000010011_0_0_00_000_000_000_0_0_00;
      patterns[2928] = 33'b1011001000010011_0_1_11_001_011_010_0_x_00;
      patterns[2929] = 33'b1011101000010011_1_1_11_001_011_010_0_x_00;
      patterns[2930] = 33'b1011101000010011_0_0_00_000_000_000_0_0_00;
      patterns[2931] = 33'b0101001000010000_0_1_xx_001_xxx_010_0_1_01;
      patterns[2932] = 33'b0101101000010000_1_1_xx_001_xxx_010_0_1_01;
      patterns[2933] = 33'b0101101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2934] = 33'b0100001000010000_0_0_xx_001_010_xxx_1_x_xx;
      patterns[2935] = 33'b0100101000010000_1_0_xx_001_010_xxx_1_x_xx;
      patterns[2936] = 33'b0100101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2937] = 33'b0000001001111100_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[2938] = 33'b0000101001111100_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[2939] = 33'b0000101001111100_0_0_00_000_000_000_0_0_00;
      patterns[2940] = 33'b1000001000010100_0_1_00_001_100_010_0_x_00;
      patterns[2941] = 33'b1000101000010100_1_1_00_001_100_010_0_x_00;
      patterns[2942] = 33'b1000101000010100_0_0_00_000_000_000_0_0_00;
      patterns[2943] = 33'b1001001000010100_0_1_01_001_100_010_0_x_00;
      patterns[2944] = 33'b1001101000010100_1_1_01_001_100_010_0_x_00;
      patterns[2945] = 33'b1001101000010100_0_0_00_000_000_000_0_0_00;
      patterns[2946] = 33'b1010001000010100_0_1_10_001_100_010_0_x_00;
      patterns[2947] = 33'b1010101000010100_1_1_10_001_100_010_0_x_00;
      patterns[2948] = 33'b1010101000010100_0_0_00_000_000_000_0_0_00;
      patterns[2949] = 33'b1011001000010100_0_1_11_001_100_010_0_x_00;
      patterns[2950] = 33'b1011101000010100_1_1_11_001_100_010_0_x_00;
      patterns[2951] = 33'b1011101000010100_0_0_00_000_000_000_0_0_00;
      patterns[2952] = 33'b0101001000010000_0_1_xx_001_xxx_010_0_1_01;
      patterns[2953] = 33'b0101101000010000_1_1_xx_001_xxx_010_0_1_01;
      patterns[2954] = 33'b0101101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2955] = 33'b0100001000010000_0_0_xx_001_010_xxx_1_x_xx;
      patterns[2956] = 33'b0100101000010000_1_0_xx_001_010_xxx_1_x_xx;
      patterns[2957] = 33'b0100101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2958] = 33'b0000001000000000_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[2959] = 33'b0000101000000000_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[2960] = 33'b0000101000000000_0_0_00_000_000_000_0_0_00;
      patterns[2961] = 33'b1000001000010101_0_1_00_001_101_010_0_x_00;
      patterns[2962] = 33'b1000101000010101_1_1_00_001_101_010_0_x_00;
      patterns[2963] = 33'b1000101000010101_0_0_00_000_000_000_0_0_00;
      patterns[2964] = 33'b1001001000010101_0_1_01_001_101_010_0_x_00;
      patterns[2965] = 33'b1001101000010101_1_1_01_001_101_010_0_x_00;
      patterns[2966] = 33'b1001101000010101_0_0_00_000_000_000_0_0_00;
      patterns[2967] = 33'b1010001000010101_0_1_10_001_101_010_0_x_00;
      patterns[2968] = 33'b1010101000010101_1_1_10_001_101_010_0_x_00;
      patterns[2969] = 33'b1010101000010101_0_0_00_000_000_000_0_0_00;
      patterns[2970] = 33'b1011001000010101_0_1_11_001_101_010_0_x_00;
      patterns[2971] = 33'b1011101000010101_1_1_11_001_101_010_0_x_00;
      patterns[2972] = 33'b1011101000010101_0_0_00_000_000_000_0_0_00;
      patterns[2973] = 33'b0101001000010000_0_1_xx_001_xxx_010_0_1_01;
      patterns[2974] = 33'b0101101000010000_1_1_xx_001_xxx_010_0_1_01;
      patterns[2975] = 33'b0101101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2976] = 33'b0100001000010000_0_0_xx_001_010_xxx_1_x_xx;
      patterns[2977] = 33'b0100101000010000_1_0_xx_001_010_xxx_1_x_xx;
      patterns[2978] = 33'b0100101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2979] = 33'b0000001011101001_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[2980] = 33'b0000101011101001_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[2981] = 33'b0000101011101001_0_0_00_000_000_000_0_0_00;
      patterns[2982] = 33'b1000001000010110_0_1_00_001_110_010_0_x_00;
      patterns[2983] = 33'b1000101000010110_1_1_00_001_110_010_0_x_00;
      patterns[2984] = 33'b1000101000010110_0_0_00_000_000_000_0_0_00;
      patterns[2985] = 33'b1001001000010110_0_1_01_001_110_010_0_x_00;
      patterns[2986] = 33'b1001101000010110_1_1_01_001_110_010_0_x_00;
      patterns[2987] = 33'b1001101000010110_0_0_00_000_000_000_0_0_00;
      patterns[2988] = 33'b1010001000010110_0_1_10_001_110_010_0_x_00;
      patterns[2989] = 33'b1010101000010110_1_1_10_001_110_010_0_x_00;
      patterns[2990] = 33'b1010101000010110_0_0_00_000_000_000_0_0_00;
      patterns[2991] = 33'b1011001000010110_0_1_11_001_110_010_0_x_00;
      patterns[2992] = 33'b1011101000010110_1_1_11_001_110_010_0_x_00;
      patterns[2993] = 33'b1011101000010110_0_0_00_000_000_000_0_0_00;
      patterns[2994] = 33'b0101001000010000_0_1_xx_001_xxx_010_0_1_01;
      patterns[2995] = 33'b0101101000010000_1_1_xx_001_xxx_010_0_1_01;
      patterns[2996] = 33'b0101101000010000_0_0_00_000_000_000_0_0_00;
      patterns[2997] = 33'b0100001000010000_0_0_xx_001_010_xxx_1_x_xx;
      patterns[2998] = 33'b0100101000010000_1_0_xx_001_010_xxx_1_x_xx;
      patterns[2999] = 33'b0100101000010000_0_0_00_000_000_000_0_0_00;
      patterns[3000] = 33'b0000001010000001_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3001] = 33'b0000101010000001_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3002] = 33'b0000101010000001_0_0_00_000_000_000_0_0_00;
      patterns[3003] = 33'b1000001000010111_0_1_00_001_111_010_0_x_00;
      patterns[3004] = 33'b1000101000010111_1_1_00_001_111_010_0_x_00;
      patterns[3005] = 33'b1000101000010111_0_0_00_000_000_000_0_0_00;
      patterns[3006] = 33'b1001001000010111_0_1_01_001_111_010_0_x_00;
      patterns[3007] = 33'b1001101000010111_1_1_01_001_111_010_0_x_00;
      patterns[3008] = 33'b1001101000010111_0_0_00_000_000_000_0_0_00;
      patterns[3009] = 33'b1010001000010111_0_1_10_001_111_010_0_x_00;
      patterns[3010] = 33'b1010101000010111_1_1_10_001_111_010_0_x_00;
      patterns[3011] = 33'b1010101000010111_0_0_00_000_000_000_0_0_00;
      patterns[3012] = 33'b1011001000010111_0_1_11_001_111_010_0_x_00;
      patterns[3013] = 33'b1011101000010111_1_1_11_001_111_010_0_x_00;
      patterns[3014] = 33'b1011101000010111_0_0_00_000_000_000_0_0_00;
      patterns[3015] = 33'b0101001000010000_0_1_xx_001_xxx_010_0_1_01;
      patterns[3016] = 33'b0101101000010000_1_1_xx_001_xxx_010_0_1_01;
      patterns[3017] = 33'b0101101000010000_0_0_00_000_000_000_0_0_00;
      patterns[3018] = 33'b0100001000010000_0_0_xx_001_010_xxx_1_x_xx;
      patterns[3019] = 33'b0100101000010000_1_0_xx_001_010_xxx_1_x_xx;
      patterns[3020] = 33'b0100101000010000_0_0_00_000_000_000_0_0_00;
      patterns[3021] = 33'b0000001011011111_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3022] = 33'b0000101011011111_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3023] = 33'b0000101011011111_0_0_00_000_000_000_0_0_00;
      patterns[3024] = 33'b1000001000100000_0_1_00_010_000_010_0_x_00;
      patterns[3025] = 33'b1000101000100000_1_1_00_010_000_010_0_x_00;
      patterns[3026] = 33'b1000101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3027] = 33'b1001001000100000_0_1_01_010_000_010_0_x_00;
      patterns[3028] = 33'b1001101000100000_1_1_01_010_000_010_0_x_00;
      patterns[3029] = 33'b1001101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3030] = 33'b1010001000100000_0_1_10_010_000_010_0_x_00;
      patterns[3031] = 33'b1010101000100000_1_1_10_010_000_010_0_x_00;
      patterns[3032] = 33'b1010101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3033] = 33'b1011001000100000_0_1_11_010_000_010_0_x_00;
      patterns[3034] = 33'b1011101000100000_1_1_11_010_000_010_0_x_00;
      patterns[3035] = 33'b1011101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3036] = 33'b0101001000100000_0_1_xx_010_xxx_010_0_1_01;
      patterns[3037] = 33'b0101101000100000_1_1_xx_010_xxx_010_0_1_01;
      patterns[3038] = 33'b0101101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3039] = 33'b0100001000100000_0_0_xx_010_010_xxx_1_x_xx;
      patterns[3040] = 33'b0100101000100000_1_0_xx_010_010_xxx_1_x_xx;
      patterns[3041] = 33'b0100101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3042] = 33'b0000001010101111_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3043] = 33'b0000101010101111_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3044] = 33'b0000101010101111_0_0_00_000_000_000_0_0_00;
      patterns[3045] = 33'b1000001000100001_0_1_00_010_001_010_0_x_00;
      patterns[3046] = 33'b1000101000100001_1_1_00_010_001_010_0_x_00;
      patterns[3047] = 33'b1000101000100001_0_0_00_000_000_000_0_0_00;
      patterns[3048] = 33'b1001001000100001_0_1_01_010_001_010_0_x_00;
      patterns[3049] = 33'b1001101000100001_1_1_01_010_001_010_0_x_00;
      patterns[3050] = 33'b1001101000100001_0_0_00_000_000_000_0_0_00;
      patterns[3051] = 33'b1010001000100001_0_1_10_010_001_010_0_x_00;
      patterns[3052] = 33'b1010101000100001_1_1_10_010_001_010_0_x_00;
      patterns[3053] = 33'b1010101000100001_0_0_00_000_000_000_0_0_00;
      patterns[3054] = 33'b1011001000100001_0_1_11_010_001_010_0_x_00;
      patterns[3055] = 33'b1011101000100001_1_1_11_010_001_010_0_x_00;
      patterns[3056] = 33'b1011101000100001_0_0_00_000_000_000_0_0_00;
      patterns[3057] = 33'b0101001000100000_0_1_xx_010_xxx_010_0_1_01;
      patterns[3058] = 33'b0101101000100000_1_1_xx_010_xxx_010_0_1_01;
      patterns[3059] = 33'b0101101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3060] = 33'b0100001000100000_0_0_xx_010_010_xxx_1_x_xx;
      patterns[3061] = 33'b0100101000100000_1_0_xx_010_010_xxx_1_x_xx;
      patterns[3062] = 33'b0100101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3063] = 33'b0000001001010100_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3064] = 33'b0000101001010100_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3065] = 33'b0000101001010100_0_0_00_000_000_000_0_0_00;
      patterns[3066] = 33'b1000001000100010_0_1_00_010_010_010_0_x_00;
      patterns[3067] = 33'b1000101000100010_1_1_00_010_010_010_0_x_00;
      patterns[3068] = 33'b1000101000100010_0_0_00_000_000_000_0_0_00;
      patterns[3069] = 33'b1001001000100010_0_1_01_010_010_010_0_x_00;
      patterns[3070] = 33'b1001101000100010_1_1_01_010_010_010_0_x_00;
      patterns[3071] = 33'b1001101000100010_0_0_00_000_000_000_0_0_00;
      patterns[3072] = 33'b1010001000100010_0_1_10_010_010_010_0_x_00;
      patterns[3073] = 33'b1010101000100010_1_1_10_010_010_010_0_x_00;
      patterns[3074] = 33'b1010101000100010_0_0_00_000_000_000_0_0_00;
      patterns[3075] = 33'b1011001000100010_0_1_11_010_010_010_0_x_00;
      patterns[3076] = 33'b1011101000100010_1_1_11_010_010_010_0_x_00;
      patterns[3077] = 33'b1011101000100010_0_0_00_000_000_000_0_0_00;
      patterns[3078] = 33'b0101001000100000_0_1_xx_010_xxx_010_0_1_01;
      patterns[3079] = 33'b0101101000100000_1_1_xx_010_xxx_010_0_1_01;
      patterns[3080] = 33'b0101101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3081] = 33'b0100001000100000_0_0_xx_010_010_xxx_1_x_xx;
      patterns[3082] = 33'b0100101000100000_1_0_xx_010_010_xxx_1_x_xx;
      patterns[3083] = 33'b0100101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3084] = 33'b0000001001000110_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3085] = 33'b0000101001000110_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3086] = 33'b0000101001000110_0_0_00_000_000_000_0_0_00;
      patterns[3087] = 33'b1000001000100011_0_1_00_010_011_010_0_x_00;
      patterns[3088] = 33'b1000101000100011_1_1_00_010_011_010_0_x_00;
      patterns[3089] = 33'b1000101000100011_0_0_00_000_000_000_0_0_00;
      patterns[3090] = 33'b1001001000100011_0_1_01_010_011_010_0_x_00;
      patterns[3091] = 33'b1001101000100011_1_1_01_010_011_010_0_x_00;
      patterns[3092] = 33'b1001101000100011_0_0_00_000_000_000_0_0_00;
      patterns[3093] = 33'b1010001000100011_0_1_10_010_011_010_0_x_00;
      patterns[3094] = 33'b1010101000100011_1_1_10_010_011_010_0_x_00;
      patterns[3095] = 33'b1010101000100011_0_0_00_000_000_000_0_0_00;
      patterns[3096] = 33'b1011001000100011_0_1_11_010_011_010_0_x_00;
      patterns[3097] = 33'b1011101000100011_1_1_11_010_011_010_0_x_00;
      patterns[3098] = 33'b1011101000100011_0_0_00_000_000_000_0_0_00;
      patterns[3099] = 33'b0101001000100000_0_1_xx_010_xxx_010_0_1_01;
      patterns[3100] = 33'b0101101000100000_1_1_xx_010_xxx_010_0_1_01;
      patterns[3101] = 33'b0101101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3102] = 33'b0100001000100000_0_0_xx_010_010_xxx_1_x_xx;
      patterns[3103] = 33'b0100101000100000_1_0_xx_010_010_xxx_1_x_xx;
      patterns[3104] = 33'b0100101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3105] = 33'b0000001000100110_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3106] = 33'b0000101000100110_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3107] = 33'b0000101000100110_0_0_00_000_000_000_0_0_00;
      patterns[3108] = 33'b1000001000100100_0_1_00_010_100_010_0_x_00;
      patterns[3109] = 33'b1000101000100100_1_1_00_010_100_010_0_x_00;
      patterns[3110] = 33'b1000101000100100_0_0_00_000_000_000_0_0_00;
      patterns[3111] = 33'b1001001000100100_0_1_01_010_100_010_0_x_00;
      patterns[3112] = 33'b1001101000100100_1_1_01_010_100_010_0_x_00;
      patterns[3113] = 33'b1001101000100100_0_0_00_000_000_000_0_0_00;
      patterns[3114] = 33'b1010001000100100_0_1_10_010_100_010_0_x_00;
      patterns[3115] = 33'b1010101000100100_1_1_10_010_100_010_0_x_00;
      patterns[3116] = 33'b1010101000100100_0_0_00_000_000_000_0_0_00;
      patterns[3117] = 33'b1011001000100100_0_1_11_010_100_010_0_x_00;
      patterns[3118] = 33'b1011101000100100_1_1_11_010_100_010_0_x_00;
      patterns[3119] = 33'b1011101000100100_0_0_00_000_000_000_0_0_00;
      patterns[3120] = 33'b0101001000100000_0_1_xx_010_xxx_010_0_1_01;
      patterns[3121] = 33'b0101101000100000_1_1_xx_010_xxx_010_0_1_01;
      patterns[3122] = 33'b0101101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3123] = 33'b0100001000100000_0_0_xx_010_010_xxx_1_x_xx;
      patterns[3124] = 33'b0100101000100000_1_0_xx_010_010_xxx_1_x_xx;
      patterns[3125] = 33'b0100101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3126] = 33'b0000001010101001_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3127] = 33'b0000101010101001_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3128] = 33'b0000101010101001_0_0_00_000_000_000_0_0_00;
      patterns[3129] = 33'b1000001000100101_0_1_00_010_101_010_0_x_00;
      patterns[3130] = 33'b1000101000100101_1_1_00_010_101_010_0_x_00;
      patterns[3131] = 33'b1000101000100101_0_0_00_000_000_000_0_0_00;
      patterns[3132] = 33'b1001001000100101_0_1_01_010_101_010_0_x_00;
      patterns[3133] = 33'b1001101000100101_1_1_01_010_101_010_0_x_00;
      patterns[3134] = 33'b1001101000100101_0_0_00_000_000_000_0_0_00;
      patterns[3135] = 33'b1010001000100101_0_1_10_010_101_010_0_x_00;
      patterns[3136] = 33'b1010101000100101_1_1_10_010_101_010_0_x_00;
      patterns[3137] = 33'b1010101000100101_0_0_00_000_000_000_0_0_00;
      patterns[3138] = 33'b1011001000100101_0_1_11_010_101_010_0_x_00;
      patterns[3139] = 33'b1011101000100101_1_1_11_010_101_010_0_x_00;
      patterns[3140] = 33'b1011101000100101_0_0_00_000_000_000_0_0_00;
      patterns[3141] = 33'b0101001000100000_0_1_xx_010_xxx_010_0_1_01;
      patterns[3142] = 33'b0101101000100000_1_1_xx_010_xxx_010_0_1_01;
      patterns[3143] = 33'b0101101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3144] = 33'b0100001000100000_0_0_xx_010_010_xxx_1_x_xx;
      patterns[3145] = 33'b0100101000100000_1_0_xx_010_010_xxx_1_x_xx;
      patterns[3146] = 33'b0100101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3147] = 33'b0000001011111010_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3148] = 33'b0000101011111010_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3149] = 33'b0000101011111010_0_0_00_000_000_000_0_0_00;
      patterns[3150] = 33'b1000001000100110_0_1_00_010_110_010_0_x_00;
      patterns[3151] = 33'b1000101000100110_1_1_00_010_110_010_0_x_00;
      patterns[3152] = 33'b1000101000100110_0_0_00_000_000_000_0_0_00;
      patterns[3153] = 33'b1001001000100110_0_1_01_010_110_010_0_x_00;
      patterns[3154] = 33'b1001101000100110_1_1_01_010_110_010_0_x_00;
      patterns[3155] = 33'b1001101000100110_0_0_00_000_000_000_0_0_00;
      patterns[3156] = 33'b1010001000100110_0_1_10_010_110_010_0_x_00;
      patterns[3157] = 33'b1010101000100110_1_1_10_010_110_010_0_x_00;
      patterns[3158] = 33'b1010101000100110_0_0_00_000_000_000_0_0_00;
      patterns[3159] = 33'b1011001000100110_0_1_11_010_110_010_0_x_00;
      patterns[3160] = 33'b1011101000100110_1_1_11_010_110_010_0_x_00;
      patterns[3161] = 33'b1011101000100110_0_0_00_000_000_000_0_0_00;
      patterns[3162] = 33'b0101001000100000_0_1_xx_010_xxx_010_0_1_01;
      patterns[3163] = 33'b0101101000100000_1_1_xx_010_xxx_010_0_1_01;
      patterns[3164] = 33'b0101101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3165] = 33'b0100001000100000_0_0_xx_010_010_xxx_1_x_xx;
      patterns[3166] = 33'b0100101000100000_1_0_xx_010_010_xxx_1_x_xx;
      patterns[3167] = 33'b0100101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3168] = 33'b0000001010101001_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3169] = 33'b0000101010101001_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3170] = 33'b0000101010101001_0_0_00_000_000_000_0_0_00;
      patterns[3171] = 33'b1000001000100111_0_1_00_010_111_010_0_x_00;
      patterns[3172] = 33'b1000101000100111_1_1_00_010_111_010_0_x_00;
      patterns[3173] = 33'b1000101000100111_0_0_00_000_000_000_0_0_00;
      patterns[3174] = 33'b1001001000100111_0_1_01_010_111_010_0_x_00;
      patterns[3175] = 33'b1001101000100111_1_1_01_010_111_010_0_x_00;
      patterns[3176] = 33'b1001101000100111_0_0_00_000_000_000_0_0_00;
      patterns[3177] = 33'b1010001000100111_0_1_10_010_111_010_0_x_00;
      patterns[3178] = 33'b1010101000100111_1_1_10_010_111_010_0_x_00;
      patterns[3179] = 33'b1010101000100111_0_0_00_000_000_000_0_0_00;
      patterns[3180] = 33'b1011001000100111_0_1_11_010_111_010_0_x_00;
      patterns[3181] = 33'b1011101000100111_1_1_11_010_111_010_0_x_00;
      patterns[3182] = 33'b1011101000100111_0_0_00_000_000_000_0_0_00;
      patterns[3183] = 33'b0101001000100000_0_1_xx_010_xxx_010_0_1_01;
      patterns[3184] = 33'b0101101000100000_1_1_xx_010_xxx_010_0_1_01;
      patterns[3185] = 33'b0101101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3186] = 33'b0100001000100000_0_0_xx_010_010_xxx_1_x_xx;
      patterns[3187] = 33'b0100101000100000_1_0_xx_010_010_xxx_1_x_xx;
      patterns[3188] = 33'b0100101000100000_0_0_00_000_000_000_0_0_00;
      patterns[3189] = 33'b0000001000000010_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3190] = 33'b0000101000000010_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3191] = 33'b0000101000000010_0_0_00_000_000_000_0_0_00;
      patterns[3192] = 33'b1000001000110000_0_1_00_011_000_010_0_x_00;
      patterns[3193] = 33'b1000101000110000_1_1_00_011_000_010_0_x_00;
      patterns[3194] = 33'b1000101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3195] = 33'b1001001000110000_0_1_01_011_000_010_0_x_00;
      patterns[3196] = 33'b1001101000110000_1_1_01_011_000_010_0_x_00;
      patterns[3197] = 33'b1001101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3198] = 33'b1010001000110000_0_1_10_011_000_010_0_x_00;
      patterns[3199] = 33'b1010101000110000_1_1_10_011_000_010_0_x_00;
      patterns[3200] = 33'b1010101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3201] = 33'b1011001000110000_0_1_11_011_000_010_0_x_00;
      patterns[3202] = 33'b1011101000110000_1_1_11_011_000_010_0_x_00;
      patterns[3203] = 33'b1011101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3204] = 33'b0101001000110000_0_1_xx_011_xxx_010_0_1_01;
      patterns[3205] = 33'b0101101000110000_1_1_xx_011_xxx_010_0_1_01;
      patterns[3206] = 33'b0101101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3207] = 33'b0100001000110000_0_0_xx_011_010_xxx_1_x_xx;
      patterns[3208] = 33'b0100101000110000_1_0_xx_011_010_xxx_1_x_xx;
      patterns[3209] = 33'b0100101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3210] = 33'b0000001000011011_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3211] = 33'b0000101000011011_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3212] = 33'b0000101000011011_0_0_00_000_000_000_0_0_00;
      patterns[3213] = 33'b1000001000110001_0_1_00_011_001_010_0_x_00;
      patterns[3214] = 33'b1000101000110001_1_1_00_011_001_010_0_x_00;
      patterns[3215] = 33'b1000101000110001_0_0_00_000_000_000_0_0_00;
      patterns[3216] = 33'b1001001000110001_0_1_01_011_001_010_0_x_00;
      patterns[3217] = 33'b1001101000110001_1_1_01_011_001_010_0_x_00;
      patterns[3218] = 33'b1001101000110001_0_0_00_000_000_000_0_0_00;
      patterns[3219] = 33'b1010001000110001_0_1_10_011_001_010_0_x_00;
      patterns[3220] = 33'b1010101000110001_1_1_10_011_001_010_0_x_00;
      patterns[3221] = 33'b1010101000110001_0_0_00_000_000_000_0_0_00;
      patterns[3222] = 33'b1011001000110001_0_1_11_011_001_010_0_x_00;
      patterns[3223] = 33'b1011101000110001_1_1_11_011_001_010_0_x_00;
      patterns[3224] = 33'b1011101000110001_0_0_00_000_000_000_0_0_00;
      patterns[3225] = 33'b0101001000110000_0_1_xx_011_xxx_010_0_1_01;
      patterns[3226] = 33'b0101101000110000_1_1_xx_011_xxx_010_0_1_01;
      patterns[3227] = 33'b0101101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3228] = 33'b0100001000110000_0_0_xx_011_010_xxx_1_x_xx;
      patterns[3229] = 33'b0100101000110000_1_0_xx_011_010_xxx_1_x_xx;
      patterns[3230] = 33'b0100101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3231] = 33'b0000001001000001_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3232] = 33'b0000101001000001_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3233] = 33'b0000101001000001_0_0_00_000_000_000_0_0_00;
      patterns[3234] = 33'b1000001000110010_0_1_00_011_010_010_0_x_00;
      patterns[3235] = 33'b1000101000110010_1_1_00_011_010_010_0_x_00;
      patterns[3236] = 33'b1000101000110010_0_0_00_000_000_000_0_0_00;
      patterns[3237] = 33'b1001001000110010_0_1_01_011_010_010_0_x_00;
      patterns[3238] = 33'b1001101000110010_1_1_01_011_010_010_0_x_00;
      patterns[3239] = 33'b1001101000110010_0_0_00_000_000_000_0_0_00;
      patterns[3240] = 33'b1010001000110010_0_1_10_011_010_010_0_x_00;
      patterns[3241] = 33'b1010101000110010_1_1_10_011_010_010_0_x_00;
      patterns[3242] = 33'b1010101000110010_0_0_00_000_000_000_0_0_00;
      patterns[3243] = 33'b1011001000110010_0_1_11_011_010_010_0_x_00;
      patterns[3244] = 33'b1011101000110010_1_1_11_011_010_010_0_x_00;
      patterns[3245] = 33'b1011101000110010_0_0_00_000_000_000_0_0_00;
      patterns[3246] = 33'b0101001000110000_0_1_xx_011_xxx_010_0_1_01;
      patterns[3247] = 33'b0101101000110000_1_1_xx_011_xxx_010_0_1_01;
      patterns[3248] = 33'b0101101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3249] = 33'b0100001000110000_0_0_xx_011_010_xxx_1_x_xx;
      patterns[3250] = 33'b0100101000110000_1_0_xx_011_010_xxx_1_x_xx;
      patterns[3251] = 33'b0100101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3252] = 33'b0000001001000001_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3253] = 33'b0000101001000001_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3254] = 33'b0000101001000001_0_0_00_000_000_000_0_0_00;
      patterns[3255] = 33'b1000001000110011_0_1_00_011_011_010_0_x_00;
      patterns[3256] = 33'b1000101000110011_1_1_00_011_011_010_0_x_00;
      patterns[3257] = 33'b1000101000110011_0_0_00_000_000_000_0_0_00;
      patterns[3258] = 33'b1001001000110011_0_1_01_011_011_010_0_x_00;
      patterns[3259] = 33'b1001101000110011_1_1_01_011_011_010_0_x_00;
      patterns[3260] = 33'b1001101000110011_0_0_00_000_000_000_0_0_00;
      patterns[3261] = 33'b1010001000110011_0_1_10_011_011_010_0_x_00;
      patterns[3262] = 33'b1010101000110011_1_1_10_011_011_010_0_x_00;
      patterns[3263] = 33'b1010101000110011_0_0_00_000_000_000_0_0_00;
      patterns[3264] = 33'b1011001000110011_0_1_11_011_011_010_0_x_00;
      patterns[3265] = 33'b1011101000110011_1_1_11_011_011_010_0_x_00;
      patterns[3266] = 33'b1011101000110011_0_0_00_000_000_000_0_0_00;
      patterns[3267] = 33'b0101001000110000_0_1_xx_011_xxx_010_0_1_01;
      patterns[3268] = 33'b0101101000110000_1_1_xx_011_xxx_010_0_1_01;
      patterns[3269] = 33'b0101101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3270] = 33'b0100001000110000_0_0_xx_011_010_xxx_1_x_xx;
      patterns[3271] = 33'b0100101000110000_1_0_xx_011_010_xxx_1_x_xx;
      patterns[3272] = 33'b0100101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3273] = 33'b0000001001010000_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3274] = 33'b0000101001010000_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3275] = 33'b0000101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3276] = 33'b1000001000110100_0_1_00_011_100_010_0_x_00;
      patterns[3277] = 33'b1000101000110100_1_1_00_011_100_010_0_x_00;
      patterns[3278] = 33'b1000101000110100_0_0_00_000_000_000_0_0_00;
      patterns[3279] = 33'b1001001000110100_0_1_01_011_100_010_0_x_00;
      patterns[3280] = 33'b1001101000110100_1_1_01_011_100_010_0_x_00;
      patterns[3281] = 33'b1001101000110100_0_0_00_000_000_000_0_0_00;
      patterns[3282] = 33'b1010001000110100_0_1_10_011_100_010_0_x_00;
      patterns[3283] = 33'b1010101000110100_1_1_10_011_100_010_0_x_00;
      patterns[3284] = 33'b1010101000110100_0_0_00_000_000_000_0_0_00;
      patterns[3285] = 33'b1011001000110100_0_1_11_011_100_010_0_x_00;
      patterns[3286] = 33'b1011101000110100_1_1_11_011_100_010_0_x_00;
      patterns[3287] = 33'b1011101000110100_0_0_00_000_000_000_0_0_00;
      patterns[3288] = 33'b0101001000110000_0_1_xx_011_xxx_010_0_1_01;
      patterns[3289] = 33'b0101101000110000_1_1_xx_011_xxx_010_0_1_01;
      patterns[3290] = 33'b0101101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3291] = 33'b0100001000110000_0_0_xx_011_010_xxx_1_x_xx;
      patterns[3292] = 33'b0100101000110000_1_0_xx_011_010_xxx_1_x_xx;
      patterns[3293] = 33'b0100101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3294] = 33'b0000001010100011_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3295] = 33'b0000101010100011_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3296] = 33'b0000101010100011_0_0_00_000_000_000_0_0_00;
      patterns[3297] = 33'b1000001000110101_0_1_00_011_101_010_0_x_00;
      patterns[3298] = 33'b1000101000110101_1_1_00_011_101_010_0_x_00;
      patterns[3299] = 33'b1000101000110101_0_0_00_000_000_000_0_0_00;
      patterns[3300] = 33'b1001001000110101_0_1_01_011_101_010_0_x_00;
      patterns[3301] = 33'b1001101000110101_1_1_01_011_101_010_0_x_00;
      patterns[3302] = 33'b1001101000110101_0_0_00_000_000_000_0_0_00;
      patterns[3303] = 33'b1010001000110101_0_1_10_011_101_010_0_x_00;
      patterns[3304] = 33'b1010101000110101_1_1_10_011_101_010_0_x_00;
      patterns[3305] = 33'b1010101000110101_0_0_00_000_000_000_0_0_00;
      patterns[3306] = 33'b1011001000110101_0_1_11_011_101_010_0_x_00;
      patterns[3307] = 33'b1011101000110101_1_1_11_011_101_010_0_x_00;
      patterns[3308] = 33'b1011101000110101_0_0_00_000_000_000_0_0_00;
      patterns[3309] = 33'b0101001000110000_0_1_xx_011_xxx_010_0_1_01;
      patterns[3310] = 33'b0101101000110000_1_1_xx_011_xxx_010_0_1_01;
      patterns[3311] = 33'b0101101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3312] = 33'b0100001000110000_0_0_xx_011_010_xxx_1_x_xx;
      patterns[3313] = 33'b0100101000110000_1_0_xx_011_010_xxx_1_x_xx;
      patterns[3314] = 33'b0100101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3315] = 33'b0000001000011010_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3316] = 33'b0000101000011010_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3317] = 33'b0000101000011010_0_0_00_000_000_000_0_0_00;
      patterns[3318] = 33'b1000001000110110_0_1_00_011_110_010_0_x_00;
      patterns[3319] = 33'b1000101000110110_1_1_00_011_110_010_0_x_00;
      patterns[3320] = 33'b1000101000110110_0_0_00_000_000_000_0_0_00;
      patterns[3321] = 33'b1001001000110110_0_1_01_011_110_010_0_x_00;
      patterns[3322] = 33'b1001101000110110_1_1_01_011_110_010_0_x_00;
      patterns[3323] = 33'b1001101000110110_0_0_00_000_000_000_0_0_00;
      patterns[3324] = 33'b1010001000110110_0_1_10_011_110_010_0_x_00;
      patterns[3325] = 33'b1010101000110110_1_1_10_011_110_010_0_x_00;
      patterns[3326] = 33'b1010101000110110_0_0_00_000_000_000_0_0_00;
      patterns[3327] = 33'b1011001000110110_0_1_11_011_110_010_0_x_00;
      patterns[3328] = 33'b1011101000110110_1_1_11_011_110_010_0_x_00;
      patterns[3329] = 33'b1011101000110110_0_0_00_000_000_000_0_0_00;
      patterns[3330] = 33'b0101001000110000_0_1_xx_011_xxx_010_0_1_01;
      patterns[3331] = 33'b0101101000110000_1_1_xx_011_xxx_010_0_1_01;
      patterns[3332] = 33'b0101101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3333] = 33'b0100001000110000_0_0_xx_011_010_xxx_1_x_xx;
      patterns[3334] = 33'b0100101000110000_1_0_xx_011_010_xxx_1_x_xx;
      patterns[3335] = 33'b0100101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3336] = 33'b0000001000010000_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3337] = 33'b0000101000010000_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3338] = 33'b0000101000010000_0_0_00_000_000_000_0_0_00;
      patterns[3339] = 33'b1000001000110111_0_1_00_011_111_010_0_x_00;
      patterns[3340] = 33'b1000101000110111_1_1_00_011_111_010_0_x_00;
      patterns[3341] = 33'b1000101000110111_0_0_00_000_000_000_0_0_00;
      patterns[3342] = 33'b1001001000110111_0_1_01_011_111_010_0_x_00;
      patterns[3343] = 33'b1001101000110111_1_1_01_011_111_010_0_x_00;
      patterns[3344] = 33'b1001101000110111_0_0_00_000_000_000_0_0_00;
      patterns[3345] = 33'b1010001000110111_0_1_10_011_111_010_0_x_00;
      patterns[3346] = 33'b1010101000110111_1_1_10_011_111_010_0_x_00;
      patterns[3347] = 33'b1010101000110111_0_0_00_000_000_000_0_0_00;
      patterns[3348] = 33'b1011001000110111_0_1_11_011_111_010_0_x_00;
      patterns[3349] = 33'b1011101000110111_1_1_11_011_111_010_0_x_00;
      patterns[3350] = 33'b1011101000110111_0_0_00_000_000_000_0_0_00;
      patterns[3351] = 33'b0101001000110000_0_1_xx_011_xxx_010_0_1_01;
      patterns[3352] = 33'b0101101000110000_1_1_xx_011_xxx_010_0_1_01;
      patterns[3353] = 33'b0101101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3354] = 33'b0100001000110000_0_0_xx_011_010_xxx_1_x_xx;
      patterns[3355] = 33'b0100101000110000_1_0_xx_011_010_xxx_1_x_xx;
      patterns[3356] = 33'b0100101000110000_0_0_00_000_000_000_0_0_00;
      patterns[3357] = 33'b0000001010000111_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3358] = 33'b0000101010000111_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3359] = 33'b0000101010000111_0_0_00_000_000_000_0_0_00;
      patterns[3360] = 33'b1000001001000000_0_1_00_100_000_010_0_x_00;
      patterns[3361] = 33'b1000101001000000_1_1_00_100_000_010_0_x_00;
      patterns[3362] = 33'b1000101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3363] = 33'b1001001001000000_0_1_01_100_000_010_0_x_00;
      patterns[3364] = 33'b1001101001000000_1_1_01_100_000_010_0_x_00;
      patterns[3365] = 33'b1001101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3366] = 33'b1010001001000000_0_1_10_100_000_010_0_x_00;
      patterns[3367] = 33'b1010101001000000_1_1_10_100_000_010_0_x_00;
      patterns[3368] = 33'b1010101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3369] = 33'b1011001001000000_0_1_11_100_000_010_0_x_00;
      patterns[3370] = 33'b1011101001000000_1_1_11_100_000_010_0_x_00;
      patterns[3371] = 33'b1011101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3372] = 33'b0101001001000000_0_1_xx_100_xxx_010_0_1_01;
      patterns[3373] = 33'b0101101001000000_1_1_xx_100_xxx_010_0_1_01;
      patterns[3374] = 33'b0101101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3375] = 33'b0100001001000000_0_0_xx_100_010_xxx_1_x_xx;
      patterns[3376] = 33'b0100101001000000_1_0_xx_100_010_xxx_1_x_xx;
      patterns[3377] = 33'b0100101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3378] = 33'b0000001010101000_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3379] = 33'b0000101010101000_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3380] = 33'b0000101010101000_0_0_00_000_000_000_0_0_00;
      patterns[3381] = 33'b1000001001000001_0_1_00_100_001_010_0_x_00;
      patterns[3382] = 33'b1000101001000001_1_1_00_100_001_010_0_x_00;
      patterns[3383] = 33'b1000101001000001_0_0_00_000_000_000_0_0_00;
      patterns[3384] = 33'b1001001001000001_0_1_01_100_001_010_0_x_00;
      patterns[3385] = 33'b1001101001000001_1_1_01_100_001_010_0_x_00;
      patterns[3386] = 33'b1001101001000001_0_0_00_000_000_000_0_0_00;
      patterns[3387] = 33'b1010001001000001_0_1_10_100_001_010_0_x_00;
      patterns[3388] = 33'b1010101001000001_1_1_10_100_001_010_0_x_00;
      patterns[3389] = 33'b1010101001000001_0_0_00_000_000_000_0_0_00;
      patterns[3390] = 33'b1011001001000001_0_1_11_100_001_010_0_x_00;
      patterns[3391] = 33'b1011101001000001_1_1_11_100_001_010_0_x_00;
      patterns[3392] = 33'b1011101001000001_0_0_00_000_000_000_0_0_00;
      patterns[3393] = 33'b0101001001000000_0_1_xx_100_xxx_010_0_1_01;
      patterns[3394] = 33'b0101101001000000_1_1_xx_100_xxx_010_0_1_01;
      patterns[3395] = 33'b0101101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3396] = 33'b0100001001000000_0_0_xx_100_010_xxx_1_x_xx;
      patterns[3397] = 33'b0100101001000000_1_0_xx_100_010_xxx_1_x_xx;
      patterns[3398] = 33'b0100101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3399] = 33'b0000001010010101_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3400] = 33'b0000101010010101_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3401] = 33'b0000101010010101_0_0_00_000_000_000_0_0_00;
      patterns[3402] = 33'b1000001001000010_0_1_00_100_010_010_0_x_00;
      patterns[3403] = 33'b1000101001000010_1_1_00_100_010_010_0_x_00;
      patterns[3404] = 33'b1000101001000010_0_0_00_000_000_000_0_0_00;
      patterns[3405] = 33'b1001001001000010_0_1_01_100_010_010_0_x_00;
      patterns[3406] = 33'b1001101001000010_1_1_01_100_010_010_0_x_00;
      patterns[3407] = 33'b1001101001000010_0_0_00_000_000_000_0_0_00;
      patterns[3408] = 33'b1010001001000010_0_1_10_100_010_010_0_x_00;
      patterns[3409] = 33'b1010101001000010_1_1_10_100_010_010_0_x_00;
      patterns[3410] = 33'b1010101001000010_0_0_00_000_000_000_0_0_00;
      patterns[3411] = 33'b1011001001000010_0_1_11_100_010_010_0_x_00;
      patterns[3412] = 33'b1011101001000010_1_1_11_100_010_010_0_x_00;
      patterns[3413] = 33'b1011101001000010_0_0_00_000_000_000_0_0_00;
      patterns[3414] = 33'b0101001001000000_0_1_xx_100_xxx_010_0_1_01;
      patterns[3415] = 33'b0101101001000000_1_1_xx_100_xxx_010_0_1_01;
      patterns[3416] = 33'b0101101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3417] = 33'b0100001001000000_0_0_xx_100_010_xxx_1_x_xx;
      patterns[3418] = 33'b0100101001000000_1_0_xx_100_010_xxx_1_x_xx;
      patterns[3419] = 33'b0100101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3420] = 33'b0000001000011111_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3421] = 33'b0000101000011111_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3422] = 33'b0000101000011111_0_0_00_000_000_000_0_0_00;
      patterns[3423] = 33'b1000001001000011_0_1_00_100_011_010_0_x_00;
      patterns[3424] = 33'b1000101001000011_1_1_00_100_011_010_0_x_00;
      patterns[3425] = 33'b1000101001000011_0_0_00_000_000_000_0_0_00;
      patterns[3426] = 33'b1001001001000011_0_1_01_100_011_010_0_x_00;
      patterns[3427] = 33'b1001101001000011_1_1_01_100_011_010_0_x_00;
      patterns[3428] = 33'b1001101001000011_0_0_00_000_000_000_0_0_00;
      patterns[3429] = 33'b1010001001000011_0_1_10_100_011_010_0_x_00;
      patterns[3430] = 33'b1010101001000011_1_1_10_100_011_010_0_x_00;
      patterns[3431] = 33'b1010101001000011_0_0_00_000_000_000_0_0_00;
      patterns[3432] = 33'b1011001001000011_0_1_11_100_011_010_0_x_00;
      patterns[3433] = 33'b1011101001000011_1_1_11_100_011_010_0_x_00;
      patterns[3434] = 33'b1011101001000011_0_0_00_000_000_000_0_0_00;
      patterns[3435] = 33'b0101001001000000_0_1_xx_100_xxx_010_0_1_01;
      patterns[3436] = 33'b0101101001000000_1_1_xx_100_xxx_010_0_1_01;
      patterns[3437] = 33'b0101101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3438] = 33'b0100001001000000_0_0_xx_100_010_xxx_1_x_xx;
      patterns[3439] = 33'b0100101001000000_1_0_xx_100_010_xxx_1_x_xx;
      patterns[3440] = 33'b0100101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3441] = 33'b0000001000010101_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3442] = 33'b0000101000010101_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3443] = 33'b0000101000010101_0_0_00_000_000_000_0_0_00;
      patterns[3444] = 33'b1000001001000100_0_1_00_100_100_010_0_x_00;
      patterns[3445] = 33'b1000101001000100_1_1_00_100_100_010_0_x_00;
      patterns[3446] = 33'b1000101001000100_0_0_00_000_000_000_0_0_00;
      patterns[3447] = 33'b1001001001000100_0_1_01_100_100_010_0_x_00;
      patterns[3448] = 33'b1001101001000100_1_1_01_100_100_010_0_x_00;
      patterns[3449] = 33'b1001101001000100_0_0_00_000_000_000_0_0_00;
      patterns[3450] = 33'b1010001001000100_0_1_10_100_100_010_0_x_00;
      patterns[3451] = 33'b1010101001000100_1_1_10_100_100_010_0_x_00;
      patterns[3452] = 33'b1010101001000100_0_0_00_000_000_000_0_0_00;
      patterns[3453] = 33'b1011001001000100_0_1_11_100_100_010_0_x_00;
      patterns[3454] = 33'b1011101001000100_1_1_11_100_100_010_0_x_00;
      patterns[3455] = 33'b1011101001000100_0_0_00_000_000_000_0_0_00;
      patterns[3456] = 33'b0101001001000000_0_1_xx_100_xxx_010_0_1_01;
      patterns[3457] = 33'b0101101001000000_1_1_xx_100_xxx_010_0_1_01;
      patterns[3458] = 33'b0101101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3459] = 33'b0100001001000000_0_0_xx_100_010_xxx_1_x_xx;
      patterns[3460] = 33'b0100101001000000_1_0_xx_100_010_xxx_1_x_xx;
      patterns[3461] = 33'b0100101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3462] = 33'b0000001001001000_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3463] = 33'b0000101001001000_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3464] = 33'b0000101001001000_0_0_00_000_000_000_0_0_00;
      patterns[3465] = 33'b1000001001000101_0_1_00_100_101_010_0_x_00;
      patterns[3466] = 33'b1000101001000101_1_1_00_100_101_010_0_x_00;
      patterns[3467] = 33'b1000101001000101_0_0_00_000_000_000_0_0_00;
      patterns[3468] = 33'b1001001001000101_0_1_01_100_101_010_0_x_00;
      patterns[3469] = 33'b1001101001000101_1_1_01_100_101_010_0_x_00;
      patterns[3470] = 33'b1001101001000101_0_0_00_000_000_000_0_0_00;
      patterns[3471] = 33'b1010001001000101_0_1_10_100_101_010_0_x_00;
      patterns[3472] = 33'b1010101001000101_1_1_10_100_101_010_0_x_00;
      patterns[3473] = 33'b1010101001000101_0_0_00_000_000_000_0_0_00;
      patterns[3474] = 33'b1011001001000101_0_1_11_100_101_010_0_x_00;
      patterns[3475] = 33'b1011101001000101_1_1_11_100_101_010_0_x_00;
      patterns[3476] = 33'b1011101001000101_0_0_00_000_000_000_0_0_00;
      patterns[3477] = 33'b0101001001000000_0_1_xx_100_xxx_010_0_1_01;
      patterns[3478] = 33'b0101101001000000_1_1_xx_100_xxx_010_0_1_01;
      patterns[3479] = 33'b0101101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3480] = 33'b0100001001000000_0_0_xx_100_010_xxx_1_x_xx;
      patterns[3481] = 33'b0100101001000000_1_0_xx_100_010_xxx_1_x_xx;
      patterns[3482] = 33'b0100101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3483] = 33'b0000001000111100_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3484] = 33'b0000101000111100_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3485] = 33'b0000101000111100_0_0_00_000_000_000_0_0_00;
      patterns[3486] = 33'b1000001001000110_0_1_00_100_110_010_0_x_00;
      patterns[3487] = 33'b1000101001000110_1_1_00_100_110_010_0_x_00;
      patterns[3488] = 33'b1000101001000110_0_0_00_000_000_000_0_0_00;
      patterns[3489] = 33'b1001001001000110_0_1_01_100_110_010_0_x_00;
      patterns[3490] = 33'b1001101001000110_1_1_01_100_110_010_0_x_00;
      patterns[3491] = 33'b1001101001000110_0_0_00_000_000_000_0_0_00;
      patterns[3492] = 33'b1010001001000110_0_1_10_100_110_010_0_x_00;
      patterns[3493] = 33'b1010101001000110_1_1_10_100_110_010_0_x_00;
      patterns[3494] = 33'b1010101001000110_0_0_00_000_000_000_0_0_00;
      patterns[3495] = 33'b1011001001000110_0_1_11_100_110_010_0_x_00;
      patterns[3496] = 33'b1011101001000110_1_1_11_100_110_010_0_x_00;
      patterns[3497] = 33'b1011101001000110_0_0_00_000_000_000_0_0_00;
      patterns[3498] = 33'b0101001001000000_0_1_xx_100_xxx_010_0_1_01;
      patterns[3499] = 33'b0101101001000000_1_1_xx_100_xxx_010_0_1_01;
      patterns[3500] = 33'b0101101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3501] = 33'b0100001001000000_0_0_xx_100_010_xxx_1_x_xx;
      patterns[3502] = 33'b0100101001000000_1_0_xx_100_010_xxx_1_x_xx;
      patterns[3503] = 33'b0100101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3504] = 33'b0000001011011010_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3505] = 33'b0000101011011010_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3506] = 33'b0000101011011010_0_0_00_000_000_000_0_0_00;
      patterns[3507] = 33'b1000001001000111_0_1_00_100_111_010_0_x_00;
      patterns[3508] = 33'b1000101001000111_1_1_00_100_111_010_0_x_00;
      patterns[3509] = 33'b1000101001000111_0_0_00_000_000_000_0_0_00;
      patterns[3510] = 33'b1001001001000111_0_1_01_100_111_010_0_x_00;
      patterns[3511] = 33'b1001101001000111_1_1_01_100_111_010_0_x_00;
      patterns[3512] = 33'b1001101001000111_0_0_00_000_000_000_0_0_00;
      patterns[3513] = 33'b1010001001000111_0_1_10_100_111_010_0_x_00;
      patterns[3514] = 33'b1010101001000111_1_1_10_100_111_010_0_x_00;
      patterns[3515] = 33'b1010101001000111_0_0_00_000_000_000_0_0_00;
      patterns[3516] = 33'b1011001001000111_0_1_11_100_111_010_0_x_00;
      patterns[3517] = 33'b1011101001000111_1_1_11_100_111_010_0_x_00;
      patterns[3518] = 33'b1011101001000111_0_0_00_000_000_000_0_0_00;
      patterns[3519] = 33'b0101001001000000_0_1_xx_100_xxx_010_0_1_01;
      patterns[3520] = 33'b0101101001000000_1_1_xx_100_xxx_010_0_1_01;
      patterns[3521] = 33'b0101101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3522] = 33'b0100001001000000_0_0_xx_100_010_xxx_1_x_xx;
      patterns[3523] = 33'b0100101001000000_1_0_xx_100_010_xxx_1_x_xx;
      patterns[3524] = 33'b0100101001000000_0_0_00_000_000_000_0_0_00;
      patterns[3525] = 33'b0000001001001000_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3526] = 33'b0000101001001000_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3527] = 33'b0000101001001000_0_0_00_000_000_000_0_0_00;
      patterns[3528] = 33'b1000001001010000_0_1_00_101_000_010_0_x_00;
      patterns[3529] = 33'b1000101001010000_1_1_00_101_000_010_0_x_00;
      patterns[3530] = 33'b1000101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3531] = 33'b1001001001010000_0_1_01_101_000_010_0_x_00;
      patterns[3532] = 33'b1001101001010000_1_1_01_101_000_010_0_x_00;
      patterns[3533] = 33'b1001101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3534] = 33'b1010001001010000_0_1_10_101_000_010_0_x_00;
      patterns[3535] = 33'b1010101001010000_1_1_10_101_000_010_0_x_00;
      patterns[3536] = 33'b1010101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3537] = 33'b1011001001010000_0_1_11_101_000_010_0_x_00;
      patterns[3538] = 33'b1011101001010000_1_1_11_101_000_010_0_x_00;
      patterns[3539] = 33'b1011101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3540] = 33'b0101001001010000_0_1_xx_101_xxx_010_0_1_01;
      patterns[3541] = 33'b0101101001010000_1_1_xx_101_xxx_010_0_1_01;
      patterns[3542] = 33'b0101101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3543] = 33'b0100001001010000_0_0_xx_101_010_xxx_1_x_xx;
      patterns[3544] = 33'b0100101001010000_1_0_xx_101_010_xxx_1_x_xx;
      patterns[3545] = 33'b0100101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3546] = 33'b0000001011101001_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3547] = 33'b0000101011101001_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3548] = 33'b0000101011101001_0_0_00_000_000_000_0_0_00;
      patterns[3549] = 33'b1000001001010001_0_1_00_101_001_010_0_x_00;
      patterns[3550] = 33'b1000101001010001_1_1_00_101_001_010_0_x_00;
      patterns[3551] = 33'b1000101001010001_0_0_00_000_000_000_0_0_00;
      patterns[3552] = 33'b1001001001010001_0_1_01_101_001_010_0_x_00;
      patterns[3553] = 33'b1001101001010001_1_1_01_101_001_010_0_x_00;
      patterns[3554] = 33'b1001101001010001_0_0_00_000_000_000_0_0_00;
      patterns[3555] = 33'b1010001001010001_0_1_10_101_001_010_0_x_00;
      patterns[3556] = 33'b1010101001010001_1_1_10_101_001_010_0_x_00;
      patterns[3557] = 33'b1010101001010001_0_0_00_000_000_000_0_0_00;
      patterns[3558] = 33'b1011001001010001_0_1_11_101_001_010_0_x_00;
      patterns[3559] = 33'b1011101001010001_1_1_11_101_001_010_0_x_00;
      patterns[3560] = 33'b1011101001010001_0_0_00_000_000_000_0_0_00;
      patterns[3561] = 33'b0101001001010000_0_1_xx_101_xxx_010_0_1_01;
      patterns[3562] = 33'b0101101001010000_1_1_xx_101_xxx_010_0_1_01;
      patterns[3563] = 33'b0101101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3564] = 33'b0100001001010000_0_0_xx_101_010_xxx_1_x_xx;
      patterns[3565] = 33'b0100101001010000_1_0_xx_101_010_xxx_1_x_xx;
      patterns[3566] = 33'b0100101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3567] = 33'b0000001010111000_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3568] = 33'b0000101010111000_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3569] = 33'b0000101010111000_0_0_00_000_000_000_0_0_00;
      patterns[3570] = 33'b1000001001010010_0_1_00_101_010_010_0_x_00;
      patterns[3571] = 33'b1000101001010010_1_1_00_101_010_010_0_x_00;
      patterns[3572] = 33'b1000101001010010_0_0_00_000_000_000_0_0_00;
      patterns[3573] = 33'b1001001001010010_0_1_01_101_010_010_0_x_00;
      patterns[3574] = 33'b1001101001010010_1_1_01_101_010_010_0_x_00;
      patterns[3575] = 33'b1001101001010010_0_0_00_000_000_000_0_0_00;
      patterns[3576] = 33'b1010001001010010_0_1_10_101_010_010_0_x_00;
      patterns[3577] = 33'b1010101001010010_1_1_10_101_010_010_0_x_00;
      patterns[3578] = 33'b1010101001010010_0_0_00_000_000_000_0_0_00;
      patterns[3579] = 33'b1011001001010010_0_1_11_101_010_010_0_x_00;
      patterns[3580] = 33'b1011101001010010_1_1_11_101_010_010_0_x_00;
      patterns[3581] = 33'b1011101001010010_0_0_00_000_000_000_0_0_00;
      patterns[3582] = 33'b0101001001010000_0_1_xx_101_xxx_010_0_1_01;
      patterns[3583] = 33'b0101101001010000_1_1_xx_101_xxx_010_0_1_01;
      patterns[3584] = 33'b0101101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3585] = 33'b0100001001010000_0_0_xx_101_010_xxx_1_x_xx;
      patterns[3586] = 33'b0100101001010000_1_0_xx_101_010_xxx_1_x_xx;
      patterns[3587] = 33'b0100101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3588] = 33'b0000001010000110_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3589] = 33'b0000101010000110_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3590] = 33'b0000101010000110_0_0_00_000_000_000_0_0_00;
      patterns[3591] = 33'b1000001001010011_0_1_00_101_011_010_0_x_00;
      patterns[3592] = 33'b1000101001010011_1_1_00_101_011_010_0_x_00;
      patterns[3593] = 33'b1000101001010011_0_0_00_000_000_000_0_0_00;
      patterns[3594] = 33'b1001001001010011_0_1_01_101_011_010_0_x_00;
      patterns[3595] = 33'b1001101001010011_1_1_01_101_011_010_0_x_00;
      patterns[3596] = 33'b1001101001010011_0_0_00_000_000_000_0_0_00;
      patterns[3597] = 33'b1010001001010011_0_1_10_101_011_010_0_x_00;
      patterns[3598] = 33'b1010101001010011_1_1_10_101_011_010_0_x_00;
      patterns[3599] = 33'b1010101001010011_0_0_00_000_000_000_0_0_00;
      patterns[3600] = 33'b1011001001010011_0_1_11_101_011_010_0_x_00;
      patterns[3601] = 33'b1011101001010011_1_1_11_101_011_010_0_x_00;
      patterns[3602] = 33'b1011101001010011_0_0_00_000_000_000_0_0_00;
      patterns[3603] = 33'b0101001001010000_0_1_xx_101_xxx_010_0_1_01;
      patterns[3604] = 33'b0101101001010000_1_1_xx_101_xxx_010_0_1_01;
      patterns[3605] = 33'b0101101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3606] = 33'b0100001001010000_0_0_xx_101_010_xxx_1_x_xx;
      patterns[3607] = 33'b0100101001010000_1_0_xx_101_010_xxx_1_x_xx;
      patterns[3608] = 33'b0100101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3609] = 33'b0000001011110001_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3610] = 33'b0000101011110001_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3611] = 33'b0000101011110001_0_0_00_000_000_000_0_0_00;
      patterns[3612] = 33'b1000001001010100_0_1_00_101_100_010_0_x_00;
      patterns[3613] = 33'b1000101001010100_1_1_00_101_100_010_0_x_00;
      patterns[3614] = 33'b1000101001010100_0_0_00_000_000_000_0_0_00;
      patterns[3615] = 33'b1001001001010100_0_1_01_101_100_010_0_x_00;
      patterns[3616] = 33'b1001101001010100_1_1_01_101_100_010_0_x_00;
      patterns[3617] = 33'b1001101001010100_0_0_00_000_000_000_0_0_00;
      patterns[3618] = 33'b1010001001010100_0_1_10_101_100_010_0_x_00;
      patterns[3619] = 33'b1010101001010100_1_1_10_101_100_010_0_x_00;
      patterns[3620] = 33'b1010101001010100_0_0_00_000_000_000_0_0_00;
      patterns[3621] = 33'b1011001001010100_0_1_11_101_100_010_0_x_00;
      patterns[3622] = 33'b1011101001010100_1_1_11_101_100_010_0_x_00;
      patterns[3623] = 33'b1011101001010100_0_0_00_000_000_000_0_0_00;
      patterns[3624] = 33'b0101001001010000_0_1_xx_101_xxx_010_0_1_01;
      patterns[3625] = 33'b0101101001010000_1_1_xx_101_xxx_010_0_1_01;
      patterns[3626] = 33'b0101101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3627] = 33'b0100001001010000_0_0_xx_101_010_xxx_1_x_xx;
      patterns[3628] = 33'b0100101001010000_1_0_xx_101_010_xxx_1_x_xx;
      patterns[3629] = 33'b0100101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3630] = 33'b0000001010100000_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3631] = 33'b0000101010100000_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3632] = 33'b0000101010100000_0_0_00_000_000_000_0_0_00;
      patterns[3633] = 33'b1000001001010101_0_1_00_101_101_010_0_x_00;
      patterns[3634] = 33'b1000101001010101_1_1_00_101_101_010_0_x_00;
      patterns[3635] = 33'b1000101001010101_0_0_00_000_000_000_0_0_00;
      patterns[3636] = 33'b1001001001010101_0_1_01_101_101_010_0_x_00;
      patterns[3637] = 33'b1001101001010101_1_1_01_101_101_010_0_x_00;
      patterns[3638] = 33'b1001101001010101_0_0_00_000_000_000_0_0_00;
      patterns[3639] = 33'b1010001001010101_0_1_10_101_101_010_0_x_00;
      patterns[3640] = 33'b1010101001010101_1_1_10_101_101_010_0_x_00;
      patterns[3641] = 33'b1010101001010101_0_0_00_000_000_000_0_0_00;
      patterns[3642] = 33'b1011001001010101_0_1_11_101_101_010_0_x_00;
      patterns[3643] = 33'b1011101001010101_1_1_11_101_101_010_0_x_00;
      patterns[3644] = 33'b1011101001010101_0_0_00_000_000_000_0_0_00;
      patterns[3645] = 33'b0101001001010000_0_1_xx_101_xxx_010_0_1_01;
      patterns[3646] = 33'b0101101001010000_1_1_xx_101_xxx_010_0_1_01;
      patterns[3647] = 33'b0101101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3648] = 33'b0100001001010000_0_0_xx_101_010_xxx_1_x_xx;
      patterns[3649] = 33'b0100101001010000_1_0_xx_101_010_xxx_1_x_xx;
      patterns[3650] = 33'b0100101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3651] = 33'b0000001010110100_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3652] = 33'b0000101010110100_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3653] = 33'b0000101010110100_0_0_00_000_000_000_0_0_00;
      patterns[3654] = 33'b1000001001010110_0_1_00_101_110_010_0_x_00;
      patterns[3655] = 33'b1000101001010110_1_1_00_101_110_010_0_x_00;
      patterns[3656] = 33'b1000101001010110_0_0_00_000_000_000_0_0_00;
      patterns[3657] = 33'b1001001001010110_0_1_01_101_110_010_0_x_00;
      patterns[3658] = 33'b1001101001010110_1_1_01_101_110_010_0_x_00;
      patterns[3659] = 33'b1001101001010110_0_0_00_000_000_000_0_0_00;
      patterns[3660] = 33'b1010001001010110_0_1_10_101_110_010_0_x_00;
      patterns[3661] = 33'b1010101001010110_1_1_10_101_110_010_0_x_00;
      patterns[3662] = 33'b1010101001010110_0_0_00_000_000_000_0_0_00;
      patterns[3663] = 33'b1011001001010110_0_1_11_101_110_010_0_x_00;
      patterns[3664] = 33'b1011101001010110_1_1_11_101_110_010_0_x_00;
      patterns[3665] = 33'b1011101001010110_0_0_00_000_000_000_0_0_00;
      patterns[3666] = 33'b0101001001010000_0_1_xx_101_xxx_010_0_1_01;
      patterns[3667] = 33'b0101101001010000_1_1_xx_101_xxx_010_0_1_01;
      patterns[3668] = 33'b0101101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3669] = 33'b0100001001010000_0_0_xx_101_010_xxx_1_x_xx;
      patterns[3670] = 33'b0100101001010000_1_0_xx_101_010_xxx_1_x_xx;
      patterns[3671] = 33'b0100101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3672] = 33'b0000001010000111_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3673] = 33'b0000101010000111_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3674] = 33'b0000101010000111_0_0_00_000_000_000_0_0_00;
      patterns[3675] = 33'b1000001001010111_0_1_00_101_111_010_0_x_00;
      patterns[3676] = 33'b1000101001010111_1_1_00_101_111_010_0_x_00;
      patterns[3677] = 33'b1000101001010111_0_0_00_000_000_000_0_0_00;
      patterns[3678] = 33'b1001001001010111_0_1_01_101_111_010_0_x_00;
      patterns[3679] = 33'b1001101001010111_1_1_01_101_111_010_0_x_00;
      patterns[3680] = 33'b1001101001010111_0_0_00_000_000_000_0_0_00;
      patterns[3681] = 33'b1010001001010111_0_1_10_101_111_010_0_x_00;
      patterns[3682] = 33'b1010101001010111_1_1_10_101_111_010_0_x_00;
      patterns[3683] = 33'b1010101001010111_0_0_00_000_000_000_0_0_00;
      patterns[3684] = 33'b1011001001010111_0_1_11_101_111_010_0_x_00;
      patterns[3685] = 33'b1011101001010111_1_1_11_101_111_010_0_x_00;
      patterns[3686] = 33'b1011101001010111_0_0_00_000_000_000_0_0_00;
      patterns[3687] = 33'b0101001001010000_0_1_xx_101_xxx_010_0_1_01;
      patterns[3688] = 33'b0101101001010000_1_1_xx_101_xxx_010_0_1_01;
      patterns[3689] = 33'b0101101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3690] = 33'b0100001001010000_0_0_xx_101_010_xxx_1_x_xx;
      patterns[3691] = 33'b0100101001010000_1_0_xx_101_010_xxx_1_x_xx;
      patterns[3692] = 33'b0100101001010000_0_0_00_000_000_000_0_0_00;
      patterns[3693] = 33'b0000001010101011_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3694] = 33'b0000101010101011_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3695] = 33'b0000101010101011_0_0_00_000_000_000_0_0_00;
      patterns[3696] = 33'b1000001001100000_0_1_00_110_000_010_0_x_00;
      patterns[3697] = 33'b1000101001100000_1_1_00_110_000_010_0_x_00;
      patterns[3698] = 33'b1000101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3699] = 33'b1001001001100000_0_1_01_110_000_010_0_x_00;
      patterns[3700] = 33'b1001101001100000_1_1_01_110_000_010_0_x_00;
      patterns[3701] = 33'b1001101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3702] = 33'b1010001001100000_0_1_10_110_000_010_0_x_00;
      patterns[3703] = 33'b1010101001100000_1_1_10_110_000_010_0_x_00;
      patterns[3704] = 33'b1010101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3705] = 33'b1011001001100000_0_1_11_110_000_010_0_x_00;
      patterns[3706] = 33'b1011101001100000_1_1_11_110_000_010_0_x_00;
      patterns[3707] = 33'b1011101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3708] = 33'b0101001001100000_0_1_xx_110_xxx_010_0_1_01;
      patterns[3709] = 33'b0101101001100000_1_1_xx_110_xxx_010_0_1_01;
      patterns[3710] = 33'b0101101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3711] = 33'b0100001001100000_0_0_xx_110_010_xxx_1_x_xx;
      patterns[3712] = 33'b0100101001100000_1_0_xx_110_010_xxx_1_x_xx;
      patterns[3713] = 33'b0100101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3714] = 33'b0000001011010110_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3715] = 33'b0000101011010110_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3716] = 33'b0000101011010110_0_0_00_000_000_000_0_0_00;
      patterns[3717] = 33'b1000001001100001_0_1_00_110_001_010_0_x_00;
      patterns[3718] = 33'b1000101001100001_1_1_00_110_001_010_0_x_00;
      patterns[3719] = 33'b1000101001100001_0_0_00_000_000_000_0_0_00;
      patterns[3720] = 33'b1001001001100001_0_1_01_110_001_010_0_x_00;
      patterns[3721] = 33'b1001101001100001_1_1_01_110_001_010_0_x_00;
      patterns[3722] = 33'b1001101001100001_0_0_00_000_000_000_0_0_00;
      patterns[3723] = 33'b1010001001100001_0_1_10_110_001_010_0_x_00;
      patterns[3724] = 33'b1010101001100001_1_1_10_110_001_010_0_x_00;
      patterns[3725] = 33'b1010101001100001_0_0_00_000_000_000_0_0_00;
      patterns[3726] = 33'b1011001001100001_0_1_11_110_001_010_0_x_00;
      patterns[3727] = 33'b1011101001100001_1_1_11_110_001_010_0_x_00;
      patterns[3728] = 33'b1011101001100001_0_0_00_000_000_000_0_0_00;
      patterns[3729] = 33'b0101001001100000_0_1_xx_110_xxx_010_0_1_01;
      patterns[3730] = 33'b0101101001100000_1_1_xx_110_xxx_010_0_1_01;
      patterns[3731] = 33'b0101101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3732] = 33'b0100001001100000_0_0_xx_110_010_xxx_1_x_xx;
      patterns[3733] = 33'b0100101001100000_1_0_xx_110_010_xxx_1_x_xx;
      patterns[3734] = 33'b0100101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3735] = 33'b0000001000001100_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3736] = 33'b0000101000001100_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3737] = 33'b0000101000001100_0_0_00_000_000_000_0_0_00;
      patterns[3738] = 33'b1000001001100010_0_1_00_110_010_010_0_x_00;
      patterns[3739] = 33'b1000101001100010_1_1_00_110_010_010_0_x_00;
      patterns[3740] = 33'b1000101001100010_0_0_00_000_000_000_0_0_00;
      patterns[3741] = 33'b1001001001100010_0_1_01_110_010_010_0_x_00;
      patterns[3742] = 33'b1001101001100010_1_1_01_110_010_010_0_x_00;
      patterns[3743] = 33'b1001101001100010_0_0_00_000_000_000_0_0_00;
      patterns[3744] = 33'b1010001001100010_0_1_10_110_010_010_0_x_00;
      patterns[3745] = 33'b1010101001100010_1_1_10_110_010_010_0_x_00;
      patterns[3746] = 33'b1010101001100010_0_0_00_000_000_000_0_0_00;
      patterns[3747] = 33'b1011001001100010_0_1_11_110_010_010_0_x_00;
      patterns[3748] = 33'b1011101001100010_1_1_11_110_010_010_0_x_00;
      patterns[3749] = 33'b1011101001100010_0_0_00_000_000_000_0_0_00;
      patterns[3750] = 33'b0101001001100000_0_1_xx_110_xxx_010_0_1_01;
      patterns[3751] = 33'b0101101001100000_1_1_xx_110_xxx_010_0_1_01;
      patterns[3752] = 33'b0101101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3753] = 33'b0100001001100000_0_0_xx_110_010_xxx_1_x_xx;
      patterns[3754] = 33'b0100101001100000_1_0_xx_110_010_xxx_1_x_xx;
      patterns[3755] = 33'b0100101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3756] = 33'b0000001010111100_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3757] = 33'b0000101010111100_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3758] = 33'b0000101010111100_0_0_00_000_000_000_0_0_00;
      patterns[3759] = 33'b1000001001100011_0_1_00_110_011_010_0_x_00;
      patterns[3760] = 33'b1000101001100011_1_1_00_110_011_010_0_x_00;
      patterns[3761] = 33'b1000101001100011_0_0_00_000_000_000_0_0_00;
      patterns[3762] = 33'b1001001001100011_0_1_01_110_011_010_0_x_00;
      patterns[3763] = 33'b1001101001100011_1_1_01_110_011_010_0_x_00;
      patterns[3764] = 33'b1001101001100011_0_0_00_000_000_000_0_0_00;
      patterns[3765] = 33'b1010001001100011_0_1_10_110_011_010_0_x_00;
      patterns[3766] = 33'b1010101001100011_1_1_10_110_011_010_0_x_00;
      patterns[3767] = 33'b1010101001100011_0_0_00_000_000_000_0_0_00;
      patterns[3768] = 33'b1011001001100011_0_1_11_110_011_010_0_x_00;
      patterns[3769] = 33'b1011101001100011_1_1_11_110_011_010_0_x_00;
      patterns[3770] = 33'b1011101001100011_0_0_00_000_000_000_0_0_00;
      patterns[3771] = 33'b0101001001100000_0_1_xx_110_xxx_010_0_1_01;
      patterns[3772] = 33'b0101101001100000_1_1_xx_110_xxx_010_0_1_01;
      patterns[3773] = 33'b0101101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3774] = 33'b0100001001100000_0_0_xx_110_010_xxx_1_x_xx;
      patterns[3775] = 33'b0100101001100000_1_0_xx_110_010_xxx_1_x_xx;
      patterns[3776] = 33'b0100101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3777] = 33'b0000001001010011_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3778] = 33'b0000101001010011_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3779] = 33'b0000101001010011_0_0_00_000_000_000_0_0_00;
      patterns[3780] = 33'b1000001001100100_0_1_00_110_100_010_0_x_00;
      patterns[3781] = 33'b1000101001100100_1_1_00_110_100_010_0_x_00;
      patterns[3782] = 33'b1000101001100100_0_0_00_000_000_000_0_0_00;
      patterns[3783] = 33'b1001001001100100_0_1_01_110_100_010_0_x_00;
      patterns[3784] = 33'b1001101001100100_1_1_01_110_100_010_0_x_00;
      patterns[3785] = 33'b1001101001100100_0_0_00_000_000_000_0_0_00;
      patterns[3786] = 33'b1010001001100100_0_1_10_110_100_010_0_x_00;
      patterns[3787] = 33'b1010101001100100_1_1_10_110_100_010_0_x_00;
      patterns[3788] = 33'b1010101001100100_0_0_00_000_000_000_0_0_00;
      patterns[3789] = 33'b1011001001100100_0_1_11_110_100_010_0_x_00;
      patterns[3790] = 33'b1011101001100100_1_1_11_110_100_010_0_x_00;
      patterns[3791] = 33'b1011101001100100_0_0_00_000_000_000_0_0_00;
      patterns[3792] = 33'b0101001001100000_0_1_xx_110_xxx_010_0_1_01;
      patterns[3793] = 33'b0101101001100000_1_1_xx_110_xxx_010_0_1_01;
      patterns[3794] = 33'b0101101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3795] = 33'b0100001001100000_0_0_xx_110_010_xxx_1_x_xx;
      patterns[3796] = 33'b0100101001100000_1_0_xx_110_010_xxx_1_x_xx;
      patterns[3797] = 33'b0100101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3798] = 33'b0000001001000111_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3799] = 33'b0000101001000111_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3800] = 33'b0000101001000111_0_0_00_000_000_000_0_0_00;
      patterns[3801] = 33'b1000001001100101_0_1_00_110_101_010_0_x_00;
      patterns[3802] = 33'b1000101001100101_1_1_00_110_101_010_0_x_00;
      patterns[3803] = 33'b1000101001100101_0_0_00_000_000_000_0_0_00;
      patterns[3804] = 33'b1001001001100101_0_1_01_110_101_010_0_x_00;
      patterns[3805] = 33'b1001101001100101_1_1_01_110_101_010_0_x_00;
      patterns[3806] = 33'b1001101001100101_0_0_00_000_000_000_0_0_00;
      patterns[3807] = 33'b1010001001100101_0_1_10_110_101_010_0_x_00;
      patterns[3808] = 33'b1010101001100101_1_1_10_110_101_010_0_x_00;
      patterns[3809] = 33'b1010101001100101_0_0_00_000_000_000_0_0_00;
      patterns[3810] = 33'b1011001001100101_0_1_11_110_101_010_0_x_00;
      patterns[3811] = 33'b1011101001100101_1_1_11_110_101_010_0_x_00;
      patterns[3812] = 33'b1011101001100101_0_0_00_000_000_000_0_0_00;
      patterns[3813] = 33'b0101001001100000_0_1_xx_110_xxx_010_0_1_01;
      patterns[3814] = 33'b0101101001100000_1_1_xx_110_xxx_010_0_1_01;
      patterns[3815] = 33'b0101101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3816] = 33'b0100001001100000_0_0_xx_110_010_xxx_1_x_xx;
      patterns[3817] = 33'b0100101001100000_1_0_xx_110_010_xxx_1_x_xx;
      patterns[3818] = 33'b0100101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3819] = 33'b0000001011011011_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3820] = 33'b0000101011011011_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3821] = 33'b0000101011011011_0_0_00_000_000_000_0_0_00;
      patterns[3822] = 33'b1000001001100110_0_1_00_110_110_010_0_x_00;
      patterns[3823] = 33'b1000101001100110_1_1_00_110_110_010_0_x_00;
      patterns[3824] = 33'b1000101001100110_0_0_00_000_000_000_0_0_00;
      patterns[3825] = 33'b1001001001100110_0_1_01_110_110_010_0_x_00;
      patterns[3826] = 33'b1001101001100110_1_1_01_110_110_010_0_x_00;
      patterns[3827] = 33'b1001101001100110_0_0_00_000_000_000_0_0_00;
      patterns[3828] = 33'b1010001001100110_0_1_10_110_110_010_0_x_00;
      patterns[3829] = 33'b1010101001100110_1_1_10_110_110_010_0_x_00;
      patterns[3830] = 33'b1010101001100110_0_0_00_000_000_000_0_0_00;
      patterns[3831] = 33'b1011001001100110_0_1_11_110_110_010_0_x_00;
      patterns[3832] = 33'b1011101001100110_1_1_11_110_110_010_0_x_00;
      patterns[3833] = 33'b1011101001100110_0_0_00_000_000_000_0_0_00;
      patterns[3834] = 33'b0101001001100000_0_1_xx_110_xxx_010_0_1_01;
      patterns[3835] = 33'b0101101001100000_1_1_xx_110_xxx_010_0_1_01;
      patterns[3836] = 33'b0101101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3837] = 33'b0100001001100000_0_0_xx_110_010_xxx_1_x_xx;
      patterns[3838] = 33'b0100101001100000_1_0_xx_110_010_xxx_1_x_xx;
      patterns[3839] = 33'b0100101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3840] = 33'b0000001000101100_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3841] = 33'b0000101000101100_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3842] = 33'b0000101000101100_0_0_00_000_000_000_0_0_00;
      patterns[3843] = 33'b1000001001100111_0_1_00_110_111_010_0_x_00;
      patterns[3844] = 33'b1000101001100111_1_1_00_110_111_010_0_x_00;
      patterns[3845] = 33'b1000101001100111_0_0_00_000_000_000_0_0_00;
      patterns[3846] = 33'b1001001001100111_0_1_01_110_111_010_0_x_00;
      patterns[3847] = 33'b1001101001100111_1_1_01_110_111_010_0_x_00;
      patterns[3848] = 33'b1001101001100111_0_0_00_000_000_000_0_0_00;
      patterns[3849] = 33'b1010001001100111_0_1_10_110_111_010_0_x_00;
      patterns[3850] = 33'b1010101001100111_1_1_10_110_111_010_0_x_00;
      patterns[3851] = 33'b1010101001100111_0_0_00_000_000_000_0_0_00;
      patterns[3852] = 33'b1011001001100111_0_1_11_110_111_010_0_x_00;
      patterns[3853] = 33'b1011101001100111_1_1_11_110_111_010_0_x_00;
      patterns[3854] = 33'b1011101001100111_0_0_00_000_000_000_0_0_00;
      patterns[3855] = 33'b0101001001100000_0_1_xx_110_xxx_010_0_1_01;
      patterns[3856] = 33'b0101101001100000_1_1_xx_110_xxx_010_0_1_01;
      patterns[3857] = 33'b0101101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3858] = 33'b0100001001100000_0_0_xx_110_010_xxx_1_x_xx;
      patterns[3859] = 33'b0100101001100000_1_0_xx_110_010_xxx_1_x_xx;
      patterns[3860] = 33'b0100101001100000_0_0_00_000_000_000_0_0_00;
      patterns[3861] = 33'b0000001011111011_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3862] = 33'b0000101011111011_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3863] = 33'b0000101011111011_0_0_00_000_000_000_0_0_00;
      patterns[3864] = 33'b1000001001110000_0_1_00_111_000_010_0_x_00;
      patterns[3865] = 33'b1000101001110000_1_1_00_111_000_010_0_x_00;
      patterns[3866] = 33'b1000101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3867] = 33'b1001001001110000_0_1_01_111_000_010_0_x_00;
      patterns[3868] = 33'b1001101001110000_1_1_01_111_000_010_0_x_00;
      patterns[3869] = 33'b1001101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3870] = 33'b1010001001110000_0_1_10_111_000_010_0_x_00;
      patterns[3871] = 33'b1010101001110000_1_1_10_111_000_010_0_x_00;
      patterns[3872] = 33'b1010101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3873] = 33'b1011001001110000_0_1_11_111_000_010_0_x_00;
      patterns[3874] = 33'b1011101001110000_1_1_11_111_000_010_0_x_00;
      patterns[3875] = 33'b1011101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3876] = 33'b0101001001110000_0_1_xx_111_xxx_010_0_1_01;
      patterns[3877] = 33'b0101101001110000_1_1_xx_111_xxx_010_0_1_01;
      patterns[3878] = 33'b0101101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3879] = 33'b0100001001110000_0_0_xx_111_010_xxx_1_x_xx;
      patterns[3880] = 33'b0100101001110000_1_0_xx_111_010_xxx_1_x_xx;
      patterns[3881] = 33'b0100101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3882] = 33'b0000001001000111_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3883] = 33'b0000101001000111_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3884] = 33'b0000101001000111_0_0_00_000_000_000_0_0_00;
      patterns[3885] = 33'b1000001001110001_0_1_00_111_001_010_0_x_00;
      patterns[3886] = 33'b1000101001110001_1_1_00_111_001_010_0_x_00;
      patterns[3887] = 33'b1000101001110001_0_0_00_000_000_000_0_0_00;
      patterns[3888] = 33'b1001001001110001_0_1_01_111_001_010_0_x_00;
      patterns[3889] = 33'b1001101001110001_1_1_01_111_001_010_0_x_00;
      patterns[3890] = 33'b1001101001110001_0_0_00_000_000_000_0_0_00;
      patterns[3891] = 33'b1010001001110001_0_1_10_111_001_010_0_x_00;
      patterns[3892] = 33'b1010101001110001_1_1_10_111_001_010_0_x_00;
      patterns[3893] = 33'b1010101001110001_0_0_00_000_000_000_0_0_00;
      patterns[3894] = 33'b1011001001110001_0_1_11_111_001_010_0_x_00;
      patterns[3895] = 33'b1011101001110001_1_1_11_111_001_010_0_x_00;
      patterns[3896] = 33'b1011101001110001_0_0_00_000_000_000_0_0_00;
      patterns[3897] = 33'b0101001001110000_0_1_xx_111_xxx_010_0_1_01;
      patterns[3898] = 33'b0101101001110000_1_1_xx_111_xxx_010_0_1_01;
      patterns[3899] = 33'b0101101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3900] = 33'b0100001001110000_0_0_xx_111_010_xxx_1_x_xx;
      patterns[3901] = 33'b0100101001110000_1_0_xx_111_010_xxx_1_x_xx;
      patterns[3902] = 33'b0100101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3903] = 33'b0000001000110100_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3904] = 33'b0000101000110100_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3905] = 33'b0000101000110100_0_0_00_000_000_000_0_0_00;
      patterns[3906] = 33'b1000001001110010_0_1_00_111_010_010_0_x_00;
      patterns[3907] = 33'b1000101001110010_1_1_00_111_010_010_0_x_00;
      patterns[3908] = 33'b1000101001110010_0_0_00_000_000_000_0_0_00;
      patterns[3909] = 33'b1001001001110010_0_1_01_111_010_010_0_x_00;
      patterns[3910] = 33'b1001101001110010_1_1_01_111_010_010_0_x_00;
      patterns[3911] = 33'b1001101001110010_0_0_00_000_000_000_0_0_00;
      patterns[3912] = 33'b1010001001110010_0_1_10_111_010_010_0_x_00;
      patterns[3913] = 33'b1010101001110010_1_1_10_111_010_010_0_x_00;
      patterns[3914] = 33'b1010101001110010_0_0_00_000_000_000_0_0_00;
      patterns[3915] = 33'b1011001001110010_0_1_11_111_010_010_0_x_00;
      patterns[3916] = 33'b1011101001110010_1_1_11_111_010_010_0_x_00;
      patterns[3917] = 33'b1011101001110010_0_0_00_000_000_000_0_0_00;
      patterns[3918] = 33'b0101001001110000_0_1_xx_111_xxx_010_0_1_01;
      patterns[3919] = 33'b0101101001110000_1_1_xx_111_xxx_010_0_1_01;
      patterns[3920] = 33'b0101101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3921] = 33'b0100001001110000_0_0_xx_111_010_xxx_1_x_xx;
      patterns[3922] = 33'b0100101001110000_1_0_xx_111_010_xxx_1_x_xx;
      patterns[3923] = 33'b0100101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3924] = 33'b0000001000111111_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3925] = 33'b0000101000111111_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3926] = 33'b0000101000111111_0_0_00_000_000_000_0_0_00;
      patterns[3927] = 33'b1000001001110011_0_1_00_111_011_010_0_x_00;
      patterns[3928] = 33'b1000101001110011_1_1_00_111_011_010_0_x_00;
      patterns[3929] = 33'b1000101001110011_0_0_00_000_000_000_0_0_00;
      patterns[3930] = 33'b1001001001110011_0_1_01_111_011_010_0_x_00;
      patterns[3931] = 33'b1001101001110011_1_1_01_111_011_010_0_x_00;
      patterns[3932] = 33'b1001101001110011_0_0_00_000_000_000_0_0_00;
      patterns[3933] = 33'b1010001001110011_0_1_10_111_011_010_0_x_00;
      patterns[3934] = 33'b1010101001110011_1_1_10_111_011_010_0_x_00;
      patterns[3935] = 33'b1010101001110011_0_0_00_000_000_000_0_0_00;
      patterns[3936] = 33'b1011001001110011_0_1_11_111_011_010_0_x_00;
      patterns[3937] = 33'b1011101001110011_1_1_11_111_011_010_0_x_00;
      patterns[3938] = 33'b1011101001110011_0_0_00_000_000_000_0_0_00;
      patterns[3939] = 33'b0101001001110000_0_1_xx_111_xxx_010_0_1_01;
      patterns[3940] = 33'b0101101001110000_1_1_xx_111_xxx_010_0_1_01;
      patterns[3941] = 33'b0101101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3942] = 33'b0100001001110000_0_0_xx_111_010_xxx_1_x_xx;
      patterns[3943] = 33'b0100101001110000_1_0_xx_111_010_xxx_1_x_xx;
      patterns[3944] = 33'b0100101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3945] = 33'b0000001001110111_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3946] = 33'b0000101001110111_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3947] = 33'b0000101001110111_0_0_00_000_000_000_0_0_00;
      patterns[3948] = 33'b1000001001110100_0_1_00_111_100_010_0_x_00;
      patterns[3949] = 33'b1000101001110100_1_1_00_111_100_010_0_x_00;
      patterns[3950] = 33'b1000101001110100_0_0_00_000_000_000_0_0_00;
      patterns[3951] = 33'b1001001001110100_0_1_01_111_100_010_0_x_00;
      patterns[3952] = 33'b1001101001110100_1_1_01_111_100_010_0_x_00;
      patterns[3953] = 33'b1001101001110100_0_0_00_000_000_000_0_0_00;
      patterns[3954] = 33'b1010001001110100_0_1_10_111_100_010_0_x_00;
      patterns[3955] = 33'b1010101001110100_1_1_10_111_100_010_0_x_00;
      patterns[3956] = 33'b1010101001110100_0_0_00_000_000_000_0_0_00;
      patterns[3957] = 33'b1011001001110100_0_1_11_111_100_010_0_x_00;
      patterns[3958] = 33'b1011101001110100_1_1_11_111_100_010_0_x_00;
      patterns[3959] = 33'b1011101001110100_0_0_00_000_000_000_0_0_00;
      patterns[3960] = 33'b0101001001110000_0_1_xx_111_xxx_010_0_1_01;
      patterns[3961] = 33'b0101101001110000_1_1_xx_111_xxx_010_0_1_01;
      patterns[3962] = 33'b0101101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3963] = 33'b0100001001110000_0_0_xx_111_010_xxx_1_x_xx;
      patterns[3964] = 33'b0100101001110000_1_0_xx_111_010_xxx_1_x_xx;
      patterns[3965] = 33'b0100101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3966] = 33'b0000001010000101_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3967] = 33'b0000101010000101_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3968] = 33'b0000101010000101_0_0_00_000_000_000_0_0_00;
      patterns[3969] = 33'b1000001001110101_0_1_00_111_101_010_0_x_00;
      patterns[3970] = 33'b1000101001110101_1_1_00_111_101_010_0_x_00;
      patterns[3971] = 33'b1000101001110101_0_0_00_000_000_000_0_0_00;
      patterns[3972] = 33'b1001001001110101_0_1_01_111_101_010_0_x_00;
      patterns[3973] = 33'b1001101001110101_1_1_01_111_101_010_0_x_00;
      patterns[3974] = 33'b1001101001110101_0_0_00_000_000_000_0_0_00;
      patterns[3975] = 33'b1010001001110101_0_1_10_111_101_010_0_x_00;
      patterns[3976] = 33'b1010101001110101_1_1_10_111_101_010_0_x_00;
      patterns[3977] = 33'b1010101001110101_0_0_00_000_000_000_0_0_00;
      patterns[3978] = 33'b1011001001110101_0_1_11_111_101_010_0_x_00;
      patterns[3979] = 33'b1011101001110101_1_1_11_111_101_010_0_x_00;
      patterns[3980] = 33'b1011101001110101_0_0_00_000_000_000_0_0_00;
      patterns[3981] = 33'b0101001001110000_0_1_xx_111_xxx_010_0_1_01;
      patterns[3982] = 33'b0101101001110000_1_1_xx_111_xxx_010_0_1_01;
      patterns[3983] = 33'b0101101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3984] = 33'b0100001001110000_0_0_xx_111_010_xxx_1_x_xx;
      patterns[3985] = 33'b0100101001110000_1_0_xx_111_010_xxx_1_x_xx;
      patterns[3986] = 33'b0100101001110000_0_0_00_000_000_000_0_0_00;
      patterns[3987] = 33'b0000001011100011_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[3988] = 33'b0000101011100011_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[3989] = 33'b0000101011100011_0_0_00_000_000_000_0_0_00;
      patterns[3990] = 33'b1000001001110110_0_1_00_111_110_010_0_x_00;
      patterns[3991] = 33'b1000101001110110_1_1_00_111_110_010_0_x_00;
      patterns[3992] = 33'b1000101001110110_0_0_00_000_000_000_0_0_00;
      patterns[3993] = 33'b1001001001110110_0_1_01_111_110_010_0_x_00;
      patterns[3994] = 33'b1001101001110110_1_1_01_111_110_010_0_x_00;
      patterns[3995] = 33'b1001101001110110_0_0_00_000_000_000_0_0_00;
      patterns[3996] = 33'b1010001001110110_0_1_10_111_110_010_0_x_00;
      patterns[3997] = 33'b1010101001110110_1_1_10_111_110_010_0_x_00;
      patterns[3998] = 33'b1010101001110110_0_0_00_000_000_000_0_0_00;
      patterns[3999] = 33'b1011001001110110_0_1_11_111_110_010_0_x_00;
      patterns[4000] = 33'b1011101001110110_1_1_11_111_110_010_0_x_00;
      patterns[4001] = 33'b1011101001110110_0_0_00_000_000_000_0_0_00;
      patterns[4002] = 33'b0101001001110000_0_1_xx_111_xxx_010_0_1_01;
      patterns[4003] = 33'b0101101001110000_1_1_xx_111_xxx_010_0_1_01;
      patterns[4004] = 33'b0101101001110000_0_0_00_000_000_000_0_0_00;
      patterns[4005] = 33'b0100001001110000_0_0_xx_111_010_xxx_1_x_xx;
      patterns[4006] = 33'b0100101001110000_1_0_xx_111_010_xxx_1_x_xx;
      patterns[4007] = 33'b0100101001110000_0_0_00_000_000_000_0_0_00;
      patterns[4008] = 33'b0000001001101000_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[4009] = 33'b0000101001101000_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[4010] = 33'b0000101001101000_0_0_00_000_000_000_0_0_00;
      patterns[4011] = 33'b1000001001110111_0_1_00_111_111_010_0_x_00;
      patterns[4012] = 33'b1000101001110111_1_1_00_111_111_010_0_x_00;
      patterns[4013] = 33'b1000101001110111_0_0_00_000_000_000_0_0_00;
      patterns[4014] = 33'b1001001001110111_0_1_01_111_111_010_0_x_00;
      patterns[4015] = 33'b1001101001110111_1_1_01_111_111_010_0_x_00;
      patterns[4016] = 33'b1001101001110111_0_0_00_000_000_000_0_0_00;
      patterns[4017] = 33'b1010001001110111_0_1_10_111_111_010_0_x_00;
      patterns[4018] = 33'b1010101001110111_1_1_10_111_111_010_0_x_00;
      patterns[4019] = 33'b1010101001110111_0_0_00_000_000_000_0_0_00;
      patterns[4020] = 33'b1011001001110111_0_1_11_111_111_010_0_x_00;
      patterns[4021] = 33'b1011101001110111_1_1_11_111_111_010_0_x_00;
      patterns[4022] = 33'b1011101001110111_0_0_00_000_000_000_0_0_00;
      patterns[4023] = 33'b0101001001110000_0_1_xx_111_xxx_010_0_1_01;
      patterns[4024] = 33'b0101101001110000_1_1_xx_111_xxx_010_0_1_01;
      patterns[4025] = 33'b0101101001110000_0_0_00_000_000_000_0_0_00;
      patterns[4026] = 33'b0100001001110000_0_0_xx_111_010_xxx_1_x_xx;
      patterns[4027] = 33'b0100101001110000_1_0_xx_111_010_xxx_1_x_xx;
      patterns[4028] = 33'b0100101001110000_0_0_00_000_000_000_0_0_00;
      patterns[4029] = 33'b0000001001000011_0_1_xx_xxx_xxx_010_0_x_10;
      patterns[4030] = 33'b0000101001000011_1_1_xx_xxx_xxx_010_0_x_10;
      patterns[4031] = 33'b0000101001000011_0_0_00_000_000_000_0_0_00;
      patterns[4032] = 33'b1000001100000000_0_1_00_000_000_011_0_x_00;
      patterns[4033] = 33'b1000101100000000_1_1_00_000_000_011_0_x_00;
      patterns[4034] = 33'b1000101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4035] = 33'b1001001100000000_0_1_01_000_000_011_0_x_00;
      patterns[4036] = 33'b1001101100000000_1_1_01_000_000_011_0_x_00;
      patterns[4037] = 33'b1001101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4038] = 33'b1010001100000000_0_1_10_000_000_011_0_x_00;
      patterns[4039] = 33'b1010101100000000_1_1_10_000_000_011_0_x_00;
      patterns[4040] = 33'b1010101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4041] = 33'b1011001100000000_0_1_11_000_000_011_0_x_00;
      patterns[4042] = 33'b1011101100000000_1_1_11_000_000_011_0_x_00;
      patterns[4043] = 33'b1011101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4044] = 33'b0101001100000000_0_1_xx_000_xxx_011_0_1_01;
      patterns[4045] = 33'b0101101100000000_1_1_xx_000_xxx_011_0_1_01;
      patterns[4046] = 33'b0101101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4047] = 33'b0100001100000000_0_0_xx_000_011_xxx_1_x_xx;
      patterns[4048] = 33'b0100101100000000_1_0_xx_000_011_xxx_1_x_xx;
      patterns[4049] = 33'b0100101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4050] = 33'b0000001111000010_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4051] = 33'b0000101111000010_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4052] = 33'b0000101111000010_0_0_00_000_000_000_0_0_00;
      patterns[4053] = 33'b1000001100000001_0_1_00_000_001_011_0_x_00;
      patterns[4054] = 33'b1000101100000001_1_1_00_000_001_011_0_x_00;
      patterns[4055] = 33'b1000101100000001_0_0_00_000_000_000_0_0_00;
      patterns[4056] = 33'b1001001100000001_0_1_01_000_001_011_0_x_00;
      patterns[4057] = 33'b1001101100000001_1_1_01_000_001_011_0_x_00;
      patterns[4058] = 33'b1001101100000001_0_0_00_000_000_000_0_0_00;
      patterns[4059] = 33'b1010001100000001_0_1_10_000_001_011_0_x_00;
      patterns[4060] = 33'b1010101100000001_1_1_10_000_001_011_0_x_00;
      patterns[4061] = 33'b1010101100000001_0_0_00_000_000_000_0_0_00;
      patterns[4062] = 33'b1011001100000001_0_1_11_000_001_011_0_x_00;
      patterns[4063] = 33'b1011101100000001_1_1_11_000_001_011_0_x_00;
      patterns[4064] = 33'b1011101100000001_0_0_00_000_000_000_0_0_00;
      patterns[4065] = 33'b0101001100000000_0_1_xx_000_xxx_011_0_1_01;
      patterns[4066] = 33'b0101101100000000_1_1_xx_000_xxx_011_0_1_01;
      patterns[4067] = 33'b0101101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4068] = 33'b0100001100000000_0_0_xx_000_011_xxx_1_x_xx;
      patterns[4069] = 33'b0100101100000000_1_0_xx_000_011_xxx_1_x_xx;
      patterns[4070] = 33'b0100101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4071] = 33'b0000001111000000_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4072] = 33'b0000101111000000_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4073] = 33'b0000101111000000_0_0_00_000_000_000_0_0_00;
      patterns[4074] = 33'b1000001100000010_0_1_00_000_010_011_0_x_00;
      patterns[4075] = 33'b1000101100000010_1_1_00_000_010_011_0_x_00;
      patterns[4076] = 33'b1000101100000010_0_0_00_000_000_000_0_0_00;
      patterns[4077] = 33'b1001001100000010_0_1_01_000_010_011_0_x_00;
      patterns[4078] = 33'b1001101100000010_1_1_01_000_010_011_0_x_00;
      patterns[4079] = 33'b1001101100000010_0_0_00_000_000_000_0_0_00;
      patterns[4080] = 33'b1010001100000010_0_1_10_000_010_011_0_x_00;
      patterns[4081] = 33'b1010101100000010_1_1_10_000_010_011_0_x_00;
      patterns[4082] = 33'b1010101100000010_0_0_00_000_000_000_0_0_00;
      patterns[4083] = 33'b1011001100000010_0_1_11_000_010_011_0_x_00;
      patterns[4084] = 33'b1011101100000010_1_1_11_000_010_011_0_x_00;
      patterns[4085] = 33'b1011101100000010_0_0_00_000_000_000_0_0_00;
      patterns[4086] = 33'b0101001100000000_0_1_xx_000_xxx_011_0_1_01;
      patterns[4087] = 33'b0101101100000000_1_1_xx_000_xxx_011_0_1_01;
      patterns[4088] = 33'b0101101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4089] = 33'b0100001100000000_0_0_xx_000_011_xxx_1_x_xx;
      patterns[4090] = 33'b0100101100000000_1_0_xx_000_011_xxx_1_x_xx;
      patterns[4091] = 33'b0100101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4092] = 33'b0000001110010101_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4093] = 33'b0000101110010101_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4094] = 33'b0000101110010101_0_0_00_000_000_000_0_0_00;
      patterns[4095] = 33'b1000001100000011_0_1_00_000_011_011_0_x_00;
      patterns[4096] = 33'b1000101100000011_1_1_00_000_011_011_0_x_00;
      patterns[4097] = 33'b1000101100000011_0_0_00_000_000_000_0_0_00;
      patterns[4098] = 33'b1001001100000011_0_1_01_000_011_011_0_x_00;
      patterns[4099] = 33'b1001101100000011_1_1_01_000_011_011_0_x_00;
      patterns[4100] = 33'b1001101100000011_0_0_00_000_000_000_0_0_00;
      patterns[4101] = 33'b1010001100000011_0_1_10_000_011_011_0_x_00;
      patterns[4102] = 33'b1010101100000011_1_1_10_000_011_011_0_x_00;
      patterns[4103] = 33'b1010101100000011_0_0_00_000_000_000_0_0_00;
      patterns[4104] = 33'b1011001100000011_0_1_11_000_011_011_0_x_00;
      patterns[4105] = 33'b1011101100000011_1_1_11_000_011_011_0_x_00;
      patterns[4106] = 33'b1011101100000011_0_0_00_000_000_000_0_0_00;
      patterns[4107] = 33'b0101001100000000_0_1_xx_000_xxx_011_0_1_01;
      patterns[4108] = 33'b0101101100000000_1_1_xx_000_xxx_011_0_1_01;
      patterns[4109] = 33'b0101101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4110] = 33'b0100001100000000_0_0_xx_000_011_xxx_1_x_xx;
      patterns[4111] = 33'b0100101100000000_1_0_xx_000_011_xxx_1_x_xx;
      patterns[4112] = 33'b0100101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4113] = 33'b0000001110001100_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4114] = 33'b0000101110001100_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4115] = 33'b0000101110001100_0_0_00_000_000_000_0_0_00;
      patterns[4116] = 33'b1000001100000100_0_1_00_000_100_011_0_x_00;
      patterns[4117] = 33'b1000101100000100_1_1_00_000_100_011_0_x_00;
      patterns[4118] = 33'b1000101100000100_0_0_00_000_000_000_0_0_00;
      patterns[4119] = 33'b1001001100000100_0_1_01_000_100_011_0_x_00;
      patterns[4120] = 33'b1001101100000100_1_1_01_000_100_011_0_x_00;
      patterns[4121] = 33'b1001101100000100_0_0_00_000_000_000_0_0_00;
      patterns[4122] = 33'b1010001100000100_0_1_10_000_100_011_0_x_00;
      patterns[4123] = 33'b1010101100000100_1_1_10_000_100_011_0_x_00;
      patterns[4124] = 33'b1010101100000100_0_0_00_000_000_000_0_0_00;
      patterns[4125] = 33'b1011001100000100_0_1_11_000_100_011_0_x_00;
      patterns[4126] = 33'b1011101100000100_1_1_11_000_100_011_0_x_00;
      patterns[4127] = 33'b1011101100000100_0_0_00_000_000_000_0_0_00;
      patterns[4128] = 33'b0101001100000000_0_1_xx_000_xxx_011_0_1_01;
      patterns[4129] = 33'b0101101100000000_1_1_xx_000_xxx_011_0_1_01;
      patterns[4130] = 33'b0101101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4131] = 33'b0100001100000000_0_0_xx_000_011_xxx_1_x_xx;
      patterns[4132] = 33'b0100101100000000_1_0_xx_000_011_xxx_1_x_xx;
      patterns[4133] = 33'b0100101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4134] = 33'b0000001111111000_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4135] = 33'b0000101111111000_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4136] = 33'b0000101111111000_0_0_00_000_000_000_0_0_00;
      patterns[4137] = 33'b1000001100000101_0_1_00_000_101_011_0_x_00;
      patterns[4138] = 33'b1000101100000101_1_1_00_000_101_011_0_x_00;
      patterns[4139] = 33'b1000101100000101_0_0_00_000_000_000_0_0_00;
      patterns[4140] = 33'b1001001100000101_0_1_01_000_101_011_0_x_00;
      patterns[4141] = 33'b1001101100000101_1_1_01_000_101_011_0_x_00;
      patterns[4142] = 33'b1001101100000101_0_0_00_000_000_000_0_0_00;
      patterns[4143] = 33'b1010001100000101_0_1_10_000_101_011_0_x_00;
      patterns[4144] = 33'b1010101100000101_1_1_10_000_101_011_0_x_00;
      patterns[4145] = 33'b1010101100000101_0_0_00_000_000_000_0_0_00;
      patterns[4146] = 33'b1011001100000101_0_1_11_000_101_011_0_x_00;
      patterns[4147] = 33'b1011101100000101_1_1_11_000_101_011_0_x_00;
      patterns[4148] = 33'b1011101100000101_0_0_00_000_000_000_0_0_00;
      patterns[4149] = 33'b0101001100000000_0_1_xx_000_xxx_011_0_1_01;
      patterns[4150] = 33'b0101101100000000_1_1_xx_000_xxx_011_0_1_01;
      patterns[4151] = 33'b0101101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4152] = 33'b0100001100000000_0_0_xx_000_011_xxx_1_x_xx;
      patterns[4153] = 33'b0100101100000000_1_0_xx_000_011_xxx_1_x_xx;
      patterns[4154] = 33'b0100101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4155] = 33'b0000001111101101_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4156] = 33'b0000101111101101_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4157] = 33'b0000101111101101_0_0_00_000_000_000_0_0_00;
      patterns[4158] = 33'b1000001100000110_0_1_00_000_110_011_0_x_00;
      patterns[4159] = 33'b1000101100000110_1_1_00_000_110_011_0_x_00;
      patterns[4160] = 33'b1000101100000110_0_0_00_000_000_000_0_0_00;
      patterns[4161] = 33'b1001001100000110_0_1_01_000_110_011_0_x_00;
      patterns[4162] = 33'b1001101100000110_1_1_01_000_110_011_0_x_00;
      patterns[4163] = 33'b1001101100000110_0_0_00_000_000_000_0_0_00;
      patterns[4164] = 33'b1010001100000110_0_1_10_000_110_011_0_x_00;
      patterns[4165] = 33'b1010101100000110_1_1_10_000_110_011_0_x_00;
      patterns[4166] = 33'b1010101100000110_0_0_00_000_000_000_0_0_00;
      patterns[4167] = 33'b1011001100000110_0_1_11_000_110_011_0_x_00;
      patterns[4168] = 33'b1011101100000110_1_1_11_000_110_011_0_x_00;
      patterns[4169] = 33'b1011101100000110_0_0_00_000_000_000_0_0_00;
      patterns[4170] = 33'b0101001100000000_0_1_xx_000_xxx_011_0_1_01;
      patterns[4171] = 33'b0101101100000000_1_1_xx_000_xxx_011_0_1_01;
      patterns[4172] = 33'b0101101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4173] = 33'b0100001100000000_0_0_xx_000_011_xxx_1_x_xx;
      patterns[4174] = 33'b0100101100000000_1_0_xx_000_011_xxx_1_x_xx;
      patterns[4175] = 33'b0100101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4176] = 33'b0000001100001110_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4177] = 33'b0000101100001110_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4178] = 33'b0000101100001110_0_0_00_000_000_000_0_0_00;
      patterns[4179] = 33'b1000001100000111_0_1_00_000_111_011_0_x_00;
      patterns[4180] = 33'b1000101100000111_1_1_00_000_111_011_0_x_00;
      patterns[4181] = 33'b1000101100000111_0_0_00_000_000_000_0_0_00;
      patterns[4182] = 33'b1001001100000111_0_1_01_000_111_011_0_x_00;
      patterns[4183] = 33'b1001101100000111_1_1_01_000_111_011_0_x_00;
      patterns[4184] = 33'b1001101100000111_0_0_00_000_000_000_0_0_00;
      patterns[4185] = 33'b1010001100000111_0_1_10_000_111_011_0_x_00;
      patterns[4186] = 33'b1010101100000111_1_1_10_000_111_011_0_x_00;
      patterns[4187] = 33'b1010101100000111_0_0_00_000_000_000_0_0_00;
      patterns[4188] = 33'b1011001100000111_0_1_11_000_111_011_0_x_00;
      patterns[4189] = 33'b1011101100000111_1_1_11_000_111_011_0_x_00;
      patterns[4190] = 33'b1011101100000111_0_0_00_000_000_000_0_0_00;
      patterns[4191] = 33'b0101001100000000_0_1_xx_000_xxx_011_0_1_01;
      patterns[4192] = 33'b0101101100000000_1_1_xx_000_xxx_011_0_1_01;
      patterns[4193] = 33'b0101101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4194] = 33'b0100001100000000_0_0_xx_000_011_xxx_1_x_xx;
      patterns[4195] = 33'b0100101100000000_1_0_xx_000_011_xxx_1_x_xx;
      patterns[4196] = 33'b0100101100000000_0_0_00_000_000_000_0_0_00;
      patterns[4197] = 33'b0000001111000111_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4198] = 33'b0000101111000111_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4199] = 33'b0000101111000111_0_0_00_000_000_000_0_0_00;
      patterns[4200] = 33'b1000001100010000_0_1_00_001_000_011_0_x_00;
      patterns[4201] = 33'b1000101100010000_1_1_00_001_000_011_0_x_00;
      patterns[4202] = 33'b1000101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4203] = 33'b1001001100010000_0_1_01_001_000_011_0_x_00;
      patterns[4204] = 33'b1001101100010000_1_1_01_001_000_011_0_x_00;
      patterns[4205] = 33'b1001101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4206] = 33'b1010001100010000_0_1_10_001_000_011_0_x_00;
      patterns[4207] = 33'b1010101100010000_1_1_10_001_000_011_0_x_00;
      patterns[4208] = 33'b1010101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4209] = 33'b1011001100010000_0_1_11_001_000_011_0_x_00;
      patterns[4210] = 33'b1011101100010000_1_1_11_001_000_011_0_x_00;
      patterns[4211] = 33'b1011101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4212] = 33'b0101001100010000_0_1_xx_001_xxx_011_0_1_01;
      patterns[4213] = 33'b0101101100010000_1_1_xx_001_xxx_011_0_1_01;
      patterns[4214] = 33'b0101101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4215] = 33'b0100001100010000_0_0_xx_001_011_xxx_1_x_xx;
      patterns[4216] = 33'b0100101100010000_1_0_xx_001_011_xxx_1_x_xx;
      patterns[4217] = 33'b0100101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4218] = 33'b0000001100100110_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4219] = 33'b0000101100100110_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4220] = 33'b0000101100100110_0_0_00_000_000_000_0_0_00;
      patterns[4221] = 33'b1000001100010001_0_1_00_001_001_011_0_x_00;
      patterns[4222] = 33'b1000101100010001_1_1_00_001_001_011_0_x_00;
      patterns[4223] = 33'b1000101100010001_0_0_00_000_000_000_0_0_00;
      patterns[4224] = 33'b1001001100010001_0_1_01_001_001_011_0_x_00;
      patterns[4225] = 33'b1001101100010001_1_1_01_001_001_011_0_x_00;
      patterns[4226] = 33'b1001101100010001_0_0_00_000_000_000_0_0_00;
      patterns[4227] = 33'b1010001100010001_0_1_10_001_001_011_0_x_00;
      patterns[4228] = 33'b1010101100010001_1_1_10_001_001_011_0_x_00;
      patterns[4229] = 33'b1010101100010001_0_0_00_000_000_000_0_0_00;
      patterns[4230] = 33'b1011001100010001_0_1_11_001_001_011_0_x_00;
      patterns[4231] = 33'b1011101100010001_1_1_11_001_001_011_0_x_00;
      patterns[4232] = 33'b1011101100010001_0_0_00_000_000_000_0_0_00;
      patterns[4233] = 33'b0101001100010000_0_1_xx_001_xxx_011_0_1_01;
      patterns[4234] = 33'b0101101100010000_1_1_xx_001_xxx_011_0_1_01;
      patterns[4235] = 33'b0101101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4236] = 33'b0100001100010000_0_0_xx_001_011_xxx_1_x_xx;
      patterns[4237] = 33'b0100101100010000_1_0_xx_001_011_xxx_1_x_xx;
      patterns[4238] = 33'b0100101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4239] = 33'b0000001101110111_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4240] = 33'b0000101101110111_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4241] = 33'b0000101101110111_0_0_00_000_000_000_0_0_00;
      patterns[4242] = 33'b1000001100010010_0_1_00_001_010_011_0_x_00;
      patterns[4243] = 33'b1000101100010010_1_1_00_001_010_011_0_x_00;
      patterns[4244] = 33'b1000101100010010_0_0_00_000_000_000_0_0_00;
      patterns[4245] = 33'b1001001100010010_0_1_01_001_010_011_0_x_00;
      patterns[4246] = 33'b1001101100010010_1_1_01_001_010_011_0_x_00;
      patterns[4247] = 33'b1001101100010010_0_0_00_000_000_000_0_0_00;
      patterns[4248] = 33'b1010001100010010_0_1_10_001_010_011_0_x_00;
      patterns[4249] = 33'b1010101100010010_1_1_10_001_010_011_0_x_00;
      patterns[4250] = 33'b1010101100010010_0_0_00_000_000_000_0_0_00;
      patterns[4251] = 33'b1011001100010010_0_1_11_001_010_011_0_x_00;
      patterns[4252] = 33'b1011101100010010_1_1_11_001_010_011_0_x_00;
      patterns[4253] = 33'b1011101100010010_0_0_00_000_000_000_0_0_00;
      patterns[4254] = 33'b0101001100010000_0_1_xx_001_xxx_011_0_1_01;
      patterns[4255] = 33'b0101101100010000_1_1_xx_001_xxx_011_0_1_01;
      patterns[4256] = 33'b0101101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4257] = 33'b0100001100010000_0_0_xx_001_011_xxx_1_x_xx;
      patterns[4258] = 33'b0100101100010000_1_0_xx_001_011_xxx_1_x_xx;
      patterns[4259] = 33'b0100101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4260] = 33'b0000001101100000_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4261] = 33'b0000101101100000_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4262] = 33'b0000101101100000_0_0_00_000_000_000_0_0_00;
      patterns[4263] = 33'b1000001100010011_0_1_00_001_011_011_0_x_00;
      patterns[4264] = 33'b1000101100010011_1_1_00_001_011_011_0_x_00;
      patterns[4265] = 33'b1000101100010011_0_0_00_000_000_000_0_0_00;
      patterns[4266] = 33'b1001001100010011_0_1_01_001_011_011_0_x_00;
      patterns[4267] = 33'b1001101100010011_1_1_01_001_011_011_0_x_00;
      patterns[4268] = 33'b1001101100010011_0_0_00_000_000_000_0_0_00;
      patterns[4269] = 33'b1010001100010011_0_1_10_001_011_011_0_x_00;
      patterns[4270] = 33'b1010101100010011_1_1_10_001_011_011_0_x_00;
      patterns[4271] = 33'b1010101100010011_0_0_00_000_000_000_0_0_00;
      patterns[4272] = 33'b1011001100010011_0_1_11_001_011_011_0_x_00;
      patterns[4273] = 33'b1011101100010011_1_1_11_001_011_011_0_x_00;
      patterns[4274] = 33'b1011101100010011_0_0_00_000_000_000_0_0_00;
      patterns[4275] = 33'b0101001100010000_0_1_xx_001_xxx_011_0_1_01;
      patterns[4276] = 33'b0101101100010000_1_1_xx_001_xxx_011_0_1_01;
      patterns[4277] = 33'b0101101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4278] = 33'b0100001100010000_0_0_xx_001_011_xxx_1_x_xx;
      patterns[4279] = 33'b0100101100010000_1_0_xx_001_011_xxx_1_x_xx;
      patterns[4280] = 33'b0100101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4281] = 33'b0000001101010110_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4282] = 33'b0000101101010110_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4283] = 33'b0000101101010110_0_0_00_000_000_000_0_0_00;
      patterns[4284] = 33'b1000001100010100_0_1_00_001_100_011_0_x_00;
      patterns[4285] = 33'b1000101100010100_1_1_00_001_100_011_0_x_00;
      patterns[4286] = 33'b1000101100010100_0_0_00_000_000_000_0_0_00;
      patterns[4287] = 33'b1001001100010100_0_1_01_001_100_011_0_x_00;
      patterns[4288] = 33'b1001101100010100_1_1_01_001_100_011_0_x_00;
      patterns[4289] = 33'b1001101100010100_0_0_00_000_000_000_0_0_00;
      patterns[4290] = 33'b1010001100010100_0_1_10_001_100_011_0_x_00;
      patterns[4291] = 33'b1010101100010100_1_1_10_001_100_011_0_x_00;
      patterns[4292] = 33'b1010101100010100_0_0_00_000_000_000_0_0_00;
      patterns[4293] = 33'b1011001100010100_0_1_11_001_100_011_0_x_00;
      patterns[4294] = 33'b1011101100010100_1_1_11_001_100_011_0_x_00;
      patterns[4295] = 33'b1011101100010100_0_0_00_000_000_000_0_0_00;
      patterns[4296] = 33'b0101001100010000_0_1_xx_001_xxx_011_0_1_01;
      patterns[4297] = 33'b0101101100010000_1_1_xx_001_xxx_011_0_1_01;
      patterns[4298] = 33'b0101101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4299] = 33'b0100001100010000_0_0_xx_001_011_xxx_1_x_xx;
      patterns[4300] = 33'b0100101100010000_1_0_xx_001_011_xxx_1_x_xx;
      patterns[4301] = 33'b0100101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4302] = 33'b0000001101111001_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4303] = 33'b0000101101111001_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4304] = 33'b0000101101111001_0_0_00_000_000_000_0_0_00;
      patterns[4305] = 33'b1000001100010101_0_1_00_001_101_011_0_x_00;
      patterns[4306] = 33'b1000101100010101_1_1_00_001_101_011_0_x_00;
      patterns[4307] = 33'b1000101100010101_0_0_00_000_000_000_0_0_00;
      patterns[4308] = 33'b1001001100010101_0_1_01_001_101_011_0_x_00;
      patterns[4309] = 33'b1001101100010101_1_1_01_001_101_011_0_x_00;
      patterns[4310] = 33'b1001101100010101_0_0_00_000_000_000_0_0_00;
      patterns[4311] = 33'b1010001100010101_0_1_10_001_101_011_0_x_00;
      patterns[4312] = 33'b1010101100010101_1_1_10_001_101_011_0_x_00;
      patterns[4313] = 33'b1010101100010101_0_0_00_000_000_000_0_0_00;
      patterns[4314] = 33'b1011001100010101_0_1_11_001_101_011_0_x_00;
      patterns[4315] = 33'b1011101100010101_1_1_11_001_101_011_0_x_00;
      patterns[4316] = 33'b1011101100010101_0_0_00_000_000_000_0_0_00;
      patterns[4317] = 33'b0101001100010000_0_1_xx_001_xxx_011_0_1_01;
      patterns[4318] = 33'b0101101100010000_1_1_xx_001_xxx_011_0_1_01;
      patterns[4319] = 33'b0101101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4320] = 33'b0100001100010000_0_0_xx_001_011_xxx_1_x_xx;
      patterns[4321] = 33'b0100101100010000_1_0_xx_001_011_xxx_1_x_xx;
      patterns[4322] = 33'b0100101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4323] = 33'b0000001110101100_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4324] = 33'b0000101110101100_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4325] = 33'b0000101110101100_0_0_00_000_000_000_0_0_00;
      patterns[4326] = 33'b1000001100010110_0_1_00_001_110_011_0_x_00;
      patterns[4327] = 33'b1000101100010110_1_1_00_001_110_011_0_x_00;
      patterns[4328] = 33'b1000101100010110_0_0_00_000_000_000_0_0_00;
      patterns[4329] = 33'b1001001100010110_0_1_01_001_110_011_0_x_00;
      patterns[4330] = 33'b1001101100010110_1_1_01_001_110_011_0_x_00;
      patterns[4331] = 33'b1001101100010110_0_0_00_000_000_000_0_0_00;
      patterns[4332] = 33'b1010001100010110_0_1_10_001_110_011_0_x_00;
      patterns[4333] = 33'b1010101100010110_1_1_10_001_110_011_0_x_00;
      patterns[4334] = 33'b1010101100010110_0_0_00_000_000_000_0_0_00;
      patterns[4335] = 33'b1011001100010110_0_1_11_001_110_011_0_x_00;
      patterns[4336] = 33'b1011101100010110_1_1_11_001_110_011_0_x_00;
      patterns[4337] = 33'b1011101100010110_0_0_00_000_000_000_0_0_00;
      patterns[4338] = 33'b0101001100010000_0_1_xx_001_xxx_011_0_1_01;
      patterns[4339] = 33'b0101101100010000_1_1_xx_001_xxx_011_0_1_01;
      patterns[4340] = 33'b0101101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4341] = 33'b0100001100010000_0_0_xx_001_011_xxx_1_x_xx;
      patterns[4342] = 33'b0100101100010000_1_0_xx_001_011_xxx_1_x_xx;
      patterns[4343] = 33'b0100101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4344] = 33'b0000001111000100_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4345] = 33'b0000101111000100_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4346] = 33'b0000101111000100_0_0_00_000_000_000_0_0_00;
      patterns[4347] = 33'b1000001100010111_0_1_00_001_111_011_0_x_00;
      patterns[4348] = 33'b1000101100010111_1_1_00_001_111_011_0_x_00;
      patterns[4349] = 33'b1000101100010111_0_0_00_000_000_000_0_0_00;
      patterns[4350] = 33'b1001001100010111_0_1_01_001_111_011_0_x_00;
      patterns[4351] = 33'b1001101100010111_1_1_01_001_111_011_0_x_00;
      patterns[4352] = 33'b1001101100010111_0_0_00_000_000_000_0_0_00;
      patterns[4353] = 33'b1010001100010111_0_1_10_001_111_011_0_x_00;
      patterns[4354] = 33'b1010101100010111_1_1_10_001_111_011_0_x_00;
      patterns[4355] = 33'b1010101100010111_0_0_00_000_000_000_0_0_00;
      patterns[4356] = 33'b1011001100010111_0_1_11_001_111_011_0_x_00;
      patterns[4357] = 33'b1011101100010111_1_1_11_001_111_011_0_x_00;
      patterns[4358] = 33'b1011101100010111_0_0_00_000_000_000_0_0_00;
      patterns[4359] = 33'b0101001100010000_0_1_xx_001_xxx_011_0_1_01;
      patterns[4360] = 33'b0101101100010000_1_1_xx_001_xxx_011_0_1_01;
      patterns[4361] = 33'b0101101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4362] = 33'b0100001100010000_0_0_xx_001_011_xxx_1_x_xx;
      patterns[4363] = 33'b0100101100010000_1_0_xx_001_011_xxx_1_x_xx;
      patterns[4364] = 33'b0100101100010000_0_0_00_000_000_000_0_0_00;
      patterns[4365] = 33'b0000001101111010_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4366] = 33'b0000101101111010_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4367] = 33'b0000101101111010_0_0_00_000_000_000_0_0_00;
      patterns[4368] = 33'b1000001100100000_0_1_00_010_000_011_0_x_00;
      patterns[4369] = 33'b1000101100100000_1_1_00_010_000_011_0_x_00;
      patterns[4370] = 33'b1000101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4371] = 33'b1001001100100000_0_1_01_010_000_011_0_x_00;
      patterns[4372] = 33'b1001101100100000_1_1_01_010_000_011_0_x_00;
      patterns[4373] = 33'b1001101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4374] = 33'b1010001100100000_0_1_10_010_000_011_0_x_00;
      patterns[4375] = 33'b1010101100100000_1_1_10_010_000_011_0_x_00;
      patterns[4376] = 33'b1010101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4377] = 33'b1011001100100000_0_1_11_010_000_011_0_x_00;
      patterns[4378] = 33'b1011101100100000_1_1_11_010_000_011_0_x_00;
      patterns[4379] = 33'b1011101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4380] = 33'b0101001100100000_0_1_xx_010_xxx_011_0_1_01;
      patterns[4381] = 33'b0101101100100000_1_1_xx_010_xxx_011_0_1_01;
      patterns[4382] = 33'b0101101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4383] = 33'b0100001100100000_0_0_xx_010_011_xxx_1_x_xx;
      patterns[4384] = 33'b0100101100100000_1_0_xx_010_011_xxx_1_x_xx;
      patterns[4385] = 33'b0100101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4386] = 33'b0000001100000101_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4387] = 33'b0000101100000101_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4388] = 33'b0000101100000101_0_0_00_000_000_000_0_0_00;
      patterns[4389] = 33'b1000001100100001_0_1_00_010_001_011_0_x_00;
      patterns[4390] = 33'b1000101100100001_1_1_00_010_001_011_0_x_00;
      patterns[4391] = 33'b1000101100100001_0_0_00_000_000_000_0_0_00;
      patterns[4392] = 33'b1001001100100001_0_1_01_010_001_011_0_x_00;
      patterns[4393] = 33'b1001101100100001_1_1_01_010_001_011_0_x_00;
      patterns[4394] = 33'b1001101100100001_0_0_00_000_000_000_0_0_00;
      patterns[4395] = 33'b1010001100100001_0_1_10_010_001_011_0_x_00;
      patterns[4396] = 33'b1010101100100001_1_1_10_010_001_011_0_x_00;
      patterns[4397] = 33'b1010101100100001_0_0_00_000_000_000_0_0_00;
      patterns[4398] = 33'b1011001100100001_0_1_11_010_001_011_0_x_00;
      patterns[4399] = 33'b1011101100100001_1_1_11_010_001_011_0_x_00;
      patterns[4400] = 33'b1011101100100001_0_0_00_000_000_000_0_0_00;
      patterns[4401] = 33'b0101001100100000_0_1_xx_010_xxx_011_0_1_01;
      patterns[4402] = 33'b0101101100100000_1_1_xx_010_xxx_011_0_1_01;
      patterns[4403] = 33'b0101101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4404] = 33'b0100001100100000_0_0_xx_010_011_xxx_1_x_xx;
      patterns[4405] = 33'b0100101100100000_1_0_xx_010_011_xxx_1_x_xx;
      patterns[4406] = 33'b0100101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4407] = 33'b0000001110111110_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4408] = 33'b0000101110111110_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4409] = 33'b0000101110111110_0_0_00_000_000_000_0_0_00;
      patterns[4410] = 33'b1000001100100010_0_1_00_010_010_011_0_x_00;
      patterns[4411] = 33'b1000101100100010_1_1_00_010_010_011_0_x_00;
      patterns[4412] = 33'b1000101100100010_0_0_00_000_000_000_0_0_00;
      patterns[4413] = 33'b1001001100100010_0_1_01_010_010_011_0_x_00;
      patterns[4414] = 33'b1001101100100010_1_1_01_010_010_011_0_x_00;
      patterns[4415] = 33'b1001101100100010_0_0_00_000_000_000_0_0_00;
      patterns[4416] = 33'b1010001100100010_0_1_10_010_010_011_0_x_00;
      patterns[4417] = 33'b1010101100100010_1_1_10_010_010_011_0_x_00;
      patterns[4418] = 33'b1010101100100010_0_0_00_000_000_000_0_0_00;
      patterns[4419] = 33'b1011001100100010_0_1_11_010_010_011_0_x_00;
      patterns[4420] = 33'b1011101100100010_1_1_11_010_010_011_0_x_00;
      patterns[4421] = 33'b1011101100100010_0_0_00_000_000_000_0_0_00;
      patterns[4422] = 33'b0101001100100000_0_1_xx_010_xxx_011_0_1_01;
      patterns[4423] = 33'b0101101100100000_1_1_xx_010_xxx_011_0_1_01;
      patterns[4424] = 33'b0101101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4425] = 33'b0100001100100000_0_0_xx_010_011_xxx_1_x_xx;
      patterns[4426] = 33'b0100101100100000_1_0_xx_010_011_xxx_1_x_xx;
      patterns[4427] = 33'b0100101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4428] = 33'b0000001100100000_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4429] = 33'b0000101100100000_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4430] = 33'b0000101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4431] = 33'b1000001100100011_0_1_00_010_011_011_0_x_00;
      patterns[4432] = 33'b1000101100100011_1_1_00_010_011_011_0_x_00;
      patterns[4433] = 33'b1000101100100011_0_0_00_000_000_000_0_0_00;
      patterns[4434] = 33'b1001001100100011_0_1_01_010_011_011_0_x_00;
      patterns[4435] = 33'b1001101100100011_1_1_01_010_011_011_0_x_00;
      patterns[4436] = 33'b1001101100100011_0_0_00_000_000_000_0_0_00;
      patterns[4437] = 33'b1010001100100011_0_1_10_010_011_011_0_x_00;
      patterns[4438] = 33'b1010101100100011_1_1_10_010_011_011_0_x_00;
      patterns[4439] = 33'b1010101100100011_0_0_00_000_000_000_0_0_00;
      patterns[4440] = 33'b1011001100100011_0_1_11_010_011_011_0_x_00;
      patterns[4441] = 33'b1011101100100011_1_1_11_010_011_011_0_x_00;
      patterns[4442] = 33'b1011101100100011_0_0_00_000_000_000_0_0_00;
      patterns[4443] = 33'b0101001100100000_0_1_xx_010_xxx_011_0_1_01;
      patterns[4444] = 33'b0101101100100000_1_1_xx_010_xxx_011_0_1_01;
      patterns[4445] = 33'b0101101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4446] = 33'b0100001100100000_0_0_xx_010_011_xxx_1_x_xx;
      patterns[4447] = 33'b0100101100100000_1_0_xx_010_011_xxx_1_x_xx;
      patterns[4448] = 33'b0100101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4449] = 33'b0000001111100100_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4450] = 33'b0000101111100100_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4451] = 33'b0000101111100100_0_0_00_000_000_000_0_0_00;
      patterns[4452] = 33'b1000001100100100_0_1_00_010_100_011_0_x_00;
      patterns[4453] = 33'b1000101100100100_1_1_00_010_100_011_0_x_00;
      patterns[4454] = 33'b1000101100100100_0_0_00_000_000_000_0_0_00;
      patterns[4455] = 33'b1001001100100100_0_1_01_010_100_011_0_x_00;
      patterns[4456] = 33'b1001101100100100_1_1_01_010_100_011_0_x_00;
      patterns[4457] = 33'b1001101100100100_0_0_00_000_000_000_0_0_00;
      patterns[4458] = 33'b1010001100100100_0_1_10_010_100_011_0_x_00;
      patterns[4459] = 33'b1010101100100100_1_1_10_010_100_011_0_x_00;
      patterns[4460] = 33'b1010101100100100_0_0_00_000_000_000_0_0_00;
      patterns[4461] = 33'b1011001100100100_0_1_11_010_100_011_0_x_00;
      patterns[4462] = 33'b1011101100100100_1_1_11_010_100_011_0_x_00;
      patterns[4463] = 33'b1011101100100100_0_0_00_000_000_000_0_0_00;
      patterns[4464] = 33'b0101001100100000_0_1_xx_010_xxx_011_0_1_01;
      patterns[4465] = 33'b0101101100100000_1_1_xx_010_xxx_011_0_1_01;
      patterns[4466] = 33'b0101101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4467] = 33'b0100001100100000_0_0_xx_010_011_xxx_1_x_xx;
      patterns[4468] = 33'b0100101100100000_1_0_xx_010_011_xxx_1_x_xx;
      patterns[4469] = 33'b0100101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4470] = 33'b0000001100100010_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4471] = 33'b0000101100100010_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4472] = 33'b0000101100100010_0_0_00_000_000_000_0_0_00;
      patterns[4473] = 33'b1000001100100101_0_1_00_010_101_011_0_x_00;
      patterns[4474] = 33'b1000101100100101_1_1_00_010_101_011_0_x_00;
      patterns[4475] = 33'b1000101100100101_0_0_00_000_000_000_0_0_00;
      patterns[4476] = 33'b1001001100100101_0_1_01_010_101_011_0_x_00;
      patterns[4477] = 33'b1001101100100101_1_1_01_010_101_011_0_x_00;
      patterns[4478] = 33'b1001101100100101_0_0_00_000_000_000_0_0_00;
      patterns[4479] = 33'b1010001100100101_0_1_10_010_101_011_0_x_00;
      patterns[4480] = 33'b1010101100100101_1_1_10_010_101_011_0_x_00;
      patterns[4481] = 33'b1010101100100101_0_0_00_000_000_000_0_0_00;
      patterns[4482] = 33'b1011001100100101_0_1_11_010_101_011_0_x_00;
      patterns[4483] = 33'b1011101100100101_1_1_11_010_101_011_0_x_00;
      patterns[4484] = 33'b1011101100100101_0_0_00_000_000_000_0_0_00;
      patterns[4485] = 33'b0101001100100000_0_1_xx_010_xxx_011_0_1_01;
      patterns[4486] = 33'b0101101100100000_1_1_xx_010_xxx_011_0_1_01;
      patterns[4487] = 33'b0101101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4488] = 33'b0100001100100000_0_0_xx_010_011_xxx_1_x_xx;
      patterns[4489] = 33'b0100101100100000_1_0_xx_010_011_xxx_1_x_xx;
      patterns[4490] = 33'b0100101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4491] = 33'b0000001100101101_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4492] = 33'b0000101100101101_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4493] = 33'b0000101100101101_0_0_00_000_000_000_0_0_00;
      patterns[4494] = 33'b1000001100100110_0_1_00_010_110_011_0_x_00;
      patterns[4495] = 33'b1000101100100110_1_1_00_010_110_011_0_x_00;
      patterns[4496] = 33'b1000101100100110_0_0_00_000_000_000_0_0_00;
      patterns[4497] = 33'b1001001100100110_0_1_01_010_110_011_0_x_00;
      patterns[4498] = 33'b1001101100100110_1_1_01_010_110_011_0_x_00;
      patterns[4499] = 33'b1001101100100110_0_0_00_000_000_000_0_0_00;
      patterns[4500] = 33'b1010001100100110_0_1_10_010_110_011_0_x_00;
      patterns[4501] = 33'b1010101100100110_1_1_10_010_110_011_0_x_00;
      patterns[4502] = 33'b1010101100100110_0_0_00_000_000_000_0_0_00;
      patterns[4503] = 33'b1011001100100110_0_1_11_010_110_011_0_x_00;
      patterns[4504] = 33'b1011101100100110_1_1_11_010_110_011_0_x_00;
      patterns[4505] = 33'b1011101100100110_0_0_00_000_000_000_0_0_00;
      patterns[4506] = 33'b0101001100100000_0_1_xx_010_xxx_011_0_1_01;
      patterns[4507] = 33'b0101101100100000_1_1_xx_010_xxx_011_0_1_01;
      patterns[4508] = 33'b0101101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4509] = 33'b0100001100100000_0_0_xx_010_011_xxx_1_x_xx;
      patterns[4510] = 33'b0100101100100000_1_0_xx_010_011_xxx_1_x_xx;
      patterns[4511] = 33'b0100101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4512] = 33'b0000001100000001_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4513] = 33'b0000101100000001_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4514] = 33'b0000101100000001_0_0_00_000_000_000_0_0_00;
      patterns[4515] = 33'b1000001100100111_0_1_00_010_111_011_0_x_00;
      patterns[4516] = 33'b1000101100100111_1_1_00_010_111_011_0_x_00;
      patterns[4517] = 33'b1000101100100111_0_0_00_000_000_000_0_0_00;
      patterns[4518] = 33'b1001001100100111_0_1_01_010_111_011_0_x_00;
      patterns[4519] = 33'b1001101100100111_1_1_01_010_111_011_0_x_00;
      patterns[4520] = 33'b1001101100100111_0_0_00_000_000_000_0_0_00;
      patterns[4521] = 33'b1010001100100111_0_1_10_010_111_011_0_x_00;
      patterns[4522] = 33'b1010101100100111_1_1_10_010_111_011_0_x_00;
      patterns[4523] = 33'b1010101100100111_0_0_00_000_000_000_0_0_00;
      patterns[4524] = 33'b1011001100100111_0_1_11_010_111_011_0_x_00;
      patterns[4525] = 33'b1011101100100111_1_1_11_010_111_011_0_x_00;
      patterns[4526] = 33'b1011101100100111_0_0_00_000_000_000_0_0_00;
      patterns[4527] = 33'b0101001100100000_0_1_xx_010_xxx_011_0_1_01;
      patterns[4528] = 33'b0101101100100000_1_1_xx_010_xxx_011_0_1_01;
      patterns[4529] = 33'b0101101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4530] = 33'b0100001100100000_0_0_xx_010_011_xxx_1_x_xx;
      patterns[4531] = 33'b0100101100100000_1_0_xx_010_011_xxx_1_x_xx;
      patterns[4532] = 33'b0100101100100000_0_0_00_000_000_000_0_0_00;
      patterns[4533] = 33'b0000001100011010_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4534] = 33'b0000101100011010_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4535] = 33'b0000101100011010_0_0_00_000_000_000_0_0_00;
      patterns[4536] = 33'b1000001100110000_0_1_00_011_000_011_0_x_00;
      patterns[4537] = 33'b1000101100110000_1_1_00_011_000_011_0_x_00;
      patterns[4538] = 33'b1000101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4539] = 33'b1001001100110000_0_1_01_011_000_011_0_x_00;
      patterns[4540] = 33'b1001101100110000_1_1_01_011_000_011_0_x_00;
      patterns[4541] = 33'b1001101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4542] = 33'b1010001100110000_0_1_10_011_000_011_0_x_00;
      patterns[4543] = 33'b1010101100110000_1_1_10_011_000_011_0_x_00;
      patterns[4544] = 33'b1010101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4545] = 33'b1011001100110000_0_1_11_011_000_011_0_x_00;
      patterns[4546] = 33'b1011101100110000_1_1_11_011_000_011_0_x_00;
      patterns[4547] = 33'b1011101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4548] = 33'b0101001100110000_0_1_xx_011_xxx_011_0_1_01;
      patterns[4549] = 33'b0101101100110000_1_1_xx_011_xxx_011_0_1_01;
      patterns[4550] = 33'b0101101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4551] = 33'b0100001100110000_0_0_xx_011_011_xxx_1_x_xx;
      patterns[4552] = 33'b0100101100110000_1_0_xx_011_011_xxx_1_x_xx;
      patterns[4553] = 33'b0100101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4554] = 33'b0000001110100111_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4555] = 33'b0000101110100111_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4556] = 33'b0000101110100111_0_0_00_000_000_000_0_0_00;
      patterns[4557] = 33'b1000001100110001_0_1_00_011_001_011_0_x_00;
      patterns[4558] = 33'b1000101100110001_1_1_00_011_001_011_0_x_00;
      patterns[4559] = 33'b1000101100110001_0_0_00_000_000_000_0_0_00;
      patterns[4560] = 33'b1001001100110001_0_1_01_011_001_011_0_x_00;
      patterns[4561] = 33'b1001101100110001_1_1_01_011_001_011_0_x_00;
      patterns[4562] = 33'b1001101100110001_0_0_00_000_000_000_0_0_00;
      patterns[4563] = 33'b1010001100110001_0_1_10_011_001_011_0_x_00;
      patterns[4564] = 33'b1010101100110001_1_1_10_011_001_011_0_x_00;
      patterns[4565] = 33'b1010101100110001_0_0_00_000_000_000_0_0_00;
      patterns[4566] = 33'b1011001100110001_0_1_11_011_001_011_0_x_00;
      patterns[4567] = 33'b1011101100110001_1_1_11_011_001_011_0_x_00;
      patterns[4568] = 33'b1011101100110001_0_0_00_000_000_000_0_0_00;
      patterns[4569] = 33'b0101001100110000_0_1_xx_011_xxx_011_0_1_01;
      patterns[4570] = 33'b0101101100110000_1_1_xx_011_xxx_011_0_1_01;
      patterns[4571] = 33'b0101101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4572] = 33'b0100001100110000_0_0_xx_011_011_xxx_1_x_xx;
      patterns[4573] = 33'b0100101100110000_1_0_xx_011_011_xxx_1_x_xx;
      patterns[4574] = 33'b0100101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4575] = 33'b0000001110110111_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4576] = 33'b0000101110110111_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4577] = 33'b0000101110110111_0_0_00_000_000_000_0_0_00;
      patterns[4578] = 33'b1000001100110010_0_1_00_011_010_011_0_x_00;
      patterns[4579] = 33'b1000101100110010_1_1_00_011_010_011_0_x_00;
      patterns[4580] = 33'b1000101100110010_0_0_00_000_000_000_0_0_00;
      patterns[4581] = 33'b1001001100110010_0_1_01_011_010_011_0_x_00;
      patterns[4582] = 33'b1001101100110010_1_1_01_011_010_011_0_x_00;
      patterns[4583] = 33'b1001101100110010_0_0_00_000_000_000_0_0_00;
      patterns[4584] = 33'b1010001100110010_0_1_10_011_010_011_0_x_00;
      patterns[4585] = 33'b1010101100110010_1_1_10_011_010_011_0_x_00;
      patterns[4586] = 33'b1010101100110010_0_0_00_000_000_000_0_0_00;
      patterns[4587] = 33'b1011001100110010_0_1_11_011_010_011_0_x_00;
      patterns[4588] = 33'b1011101100110010_1_1_11_011_010_011_0_x_00;
      patterns[4589] = 33'b1011101100110010_0_0_00_000_000_000_0_0_00;
      patterns[4590] = 33'b0101001100110000_0_1_xx_011_xxx_011_0_1_01;
      patterns[4591] = 33'b0101101100110000_1_1_xx_011_xxx_011_0_1_01;
      patterns[4592] = 33'b0101101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4593] = 33'b0100001100110000_0_0_xx_011_011_xxx_1_x_xx;
      patterns[4594] = 33'b0100101100110000_1_0_xx_011_011_xxx_1_x_xx;
      patterns[4595] = 33'b0100101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4596] = 33'b0000001100101000_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4597] = 33'b0000101100101000_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4598] = 33'b0000101100101000_0_0_00_000_000_000_0_0_00;
      patterns[4599] = 33'b1000001100110011_0_1_00_011_011_011_0_x_00;
      patterns[4600] = 33'b1000101100110011_1_1_00_011_011_011_0_x_00;
      patterns[4601] = 33'b1000101100110011_0_0_00_000_000_000_0_0_00;
      patterns[4602] = 33'b1001001100110011_0_1_01_011_011_011_0_x_00;
      patterns[4603] = 33'b1001101100110011_1_1_01_011_011_011_0_x_00;
      patterns[4604] = 33'b1001101100110011_0_0_00_000_000_000_0_0_00;
      patterns[4605] = 33'b1010001100110011_0_1_10_011_011_011_0_x_00;
      patterns[4606] = 33'b1010101100110011_1_1_10_011_011_011_0_x_00;
      patterns[4607] = 33'b1010101100110011_0_0_00_000_000_000_0_0_00;
      patterns[4608] = 33'b1011001100110011_0_1_11_011_011_011_0_x_00;
      patterns[4609] = 33'b1011101100110011_1_1_11_011_011_011_0_x_00;
      patterns[4610] = 33'b1011101100110011_0_0_00_000_000_000_0_0_00;
      patterns[4611] = 33'b0101001100110000_0_1_xx_011_xxx_011_0_1_01;
      patterns[4612] = 33'b0101101100110000_1_1_xx_011_xxx_011_0_1_01;
      patterns[4613] = 33'b0101101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4614] = 33'b0100001100110000_0_0_xx_011_011_xxx_1_x_xx;
      patterns[4615] = 33'b0100101100110000_1_0_xx_011_011_xxx_1_x_xx;
      patterns[4616] = 33'b0100101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4617] = 33'b0000001100000010_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4618] = 33'b0000101100000010_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4619] = 33'b0000101100000010_0_0_00_000_000_000_0_0_00;
      patterns[4620] = 33'b1000001100110100_0_1_00_011_100_011_0_x_00;
      patterns[4621] = 33'b1000101100110100_1_1_00_011_100_011_0_x_00;
      patterns[4622] = 33'b1000101100110100_0_0_00_000_000_000_0_0_00;
      patterns[4623] = 33'b1001001100110100_0_1_01_011_100_011_0_x_00;
      patterns[4624] = 33'b1001101100110100_1_1_01_011_100_011_0_x_00;
      patterns[4625] = 33'b1001101100110100_0_0_00_000_000_000_0_0_00;
      patterns[4626] = 33'b1010001100110100_0_1_10_011_100_011_0_x_00;
      patterns[4627] = 33'b1010101100110100_1_1_10_011_100_011_0_x_00;
      patterns[4628] = 33'b1010101100110100_0_0_00_000_000_000_0_0_00;
      patterns[4629] = 33'b1011001100110100_0_1_11_011_100_011_0_x_00;
      patterns[4630] = 33'b1011101100110100_1_1_11_011_100_011_0_x_00;
      patterns[4631] = 33'b1011101100110100_0_0_00_000_000_000_0_0_00;
      patterns[4632] = 33'b0101001100110000_0_1_xx_011_xxx_011_0_1_01;
      patterns[4633] = 33'b0101101100110000_1_1_xx_011_xxx_011_0_1_01;
      patterns[4634] = 33'b0101101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4635] = 33'b0100001100110000_0_0_xx_011_011_xxx_1_x_xx;
      patterns[4636] = 33'b0100101100110000_1_0_xx_011_011_xxx_1_x_xx;
      patterns[4637] = 33'b0100101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4638] = 33'b0000001110100111_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4639] = 33'b0000101110100111_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4640] = 33'b0000101110100111_0_0_00_000_000_000_0_0_00;
      patterns[4641] = 33'b1000001100110101_0_1_00_011_101_011_0_x_00;
      patterns[4642] = 33'b1000101100110101_1_1_00_011_101_011_0_x_00;
      patterns[4643] = 33'b1000101100110101_0_0_00_000_000_000_0_0_00;
      patterns[4644] = 33'b1001001100110101_0_1_01_011_101_011_0_x_00;
      patterns[4645] = 33'b1001101100110101_1_1_01_011_101_011_0_x_00;
      patterns[4646] = 33'b1001101100110101_0_0_00_000_000_000_0_0_00;
      patterns[4647] = 33'b1010001100110101_0_1_10_011_101_011_0_x_00;
      patterns[4648] = 33'b1010101100110101_1_1_10_011_101_011_0_x_00;
      patterns[4649] = 33'b1010101100110101_0_0_00_000_000_000_0_0_00;
      patterns[4650] = 33'b1011001100110101_0_1_11_011_101_011_0_x_00;
      patterns[4651] = 33'b1011101100110101_1_1_11_011_101_011_0_x_00;
      patterns[4652] = 33'b1011101100110101_0_0_00_000_000_000_0_0_00;
      patterns[4653] = 33'b0101001100110000_0_1_xx_011_xxx_011_0_1_01;
      patterns[4654] = 33'b0101101100110000_1_1_xx_011_xxx_011_0_1_01;
      patterns[4655] = 33'b0101101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4656] = 33'b0100001100110000_0_0_xx_011_011_xxx_1_x_xx;
      patterns[4657] = 33'b0100101100110000_1_0_xx_011_011_xxx_1_x_xx;
      patterns[4658] = 33'b0100101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4659] = 33'b0000001110010100_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4660] = 33'b0000101110010100_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4661] = 33'b0000101110010100_0_0_00_000_000_000_0_0_00;
      patterns[4662] = 33'b1000001100110110_0_1_00_011_110_011_0_x_00;
      patterns[4663] = 33'b1000101100110110_1_1_00_011_110_011_0_x_00;
      patterns[4664] = 33'b1000101100110110_0_0_00_000_000_000_0_0_00;
      patterns[4665] = 33'b1001001100110110_0_1_01_011_110_011_0_x_00;
      patterns[4666] = 33'b1001101100110110_1_1_01_011_110_011_0_x_00;
      patterns[4667] = 33'b1001101100110110_0_0_00_000_000_000_0_0_00;
      patterns[4668] = 33'b1010001100110110_0_1_10_011_110_011_0_x_00;
      patterns[4669] = 33'b1010101100110110_1_1_10_011_110_011_0_x_00;
      patterns[4670] = 33'b1010101100110110_0_0_00_000_000_000_0_0_00;
      patterns[4671] = 33'b1011001100110110_0_1_11_011_110_011_0_x_00;
      patterns[4672] = 33'b1011101100110110_1_1_11_011_110_011_0_x_00;
      patterns[4673] = 33'b1011101100110110_0_0_00_000_000_000_0_0_00;
      patterns[4674] = 33'b0101001100110000_0_1_xx_011_xxx_011_0_1_01;
      patterns[4675] = 33'b0101101100110000_1_1_xx_011_xxx_011_0_1_01;
      patterns[4676] = 33'b0101101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4677] = 33'b0100001100110000_0_0_xx_011_011_xxx_1_x_xx;
      patterns[4678] = 33'b0100101100110000_1_0_xx_011_011_xxx_1_x_xx;
      patterns[4679] = 33'b0100101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4680] = 33'b0000001100110111_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4681] = 33'b0000101100110111_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4682] = 33'b0000101100110111_0_0_00_000_000_000_0_0_00;
      patterns[4683] = 33'b1000001100110111_0_1_00_011_111_011_0_x_00;
      patterns[4684] = 33'b1000101100110111_1_1_00_011_111_011_0_x_00;
      patterns[4685] = 33'b1000101100110111_0_0_00_000_000_000_0_0_00;
      patterns[4686] = 33'b1001001100110111_0_1_01_011_111_011_0_x_00;
      patterns[4687] = 33'b1001101100110111_1_1_01_011_111_011_0_x_00;
      patterns[4688] = 33'b1001101100110111_0_0_00_000_000_000_0_0_00;
      patterns[4689] = 33'b1010001100110111_0_1_10_011_111_011_0_x_00;
      patterns[4690] = 33'b1010101100110111_1_1_10_011_111_011_0_x_00;
      patterns[4691] = 33'b1010101100110111_0_0_00_000_000_000_0_0_00;
      patterns[4692] = 33'b1011001100110111_0_1_11_011_111_011_0_x_00;
      patterns[4693] = 33'b1011101100110111_1_1_11_011_111_011_0_x_00;
      patterns[4694] = 33'b1011101100110111_0_0_00_000_000_000_0_0_00;
      patterns[4695] = 33'b0101001100110000_0_1_xx_011_xxx_011_0_1_01;
      patterns[4696] = 33'b0101101100110000_1_1_xx_011_xxx_011_0_1_01;
      patterns[4697] = 33'b0101101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4698] = 33'b0100001100110000_0_0_xx_011_011_xxx_1_x_xx;
      patterns[4699] = 33'b0100101100110000_1_0_xx_011_011_xxx_1_x_xx;
      patterns[4700] = 33'b0100101100110000_0_0_00_000_000_000_0_0_00;
      patterns[4701] = 33'b0000001111000100_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4702] = 33'b0000101111000100_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4703] = 33'b0000101111000100_0_0_00_000_000_000_0_0_00;
      patterns[4704] = 33'b1000001101000000_0_1_00_100_000_011_0_x_00;
      patterns[4705] = 33'b1000101101000000_1_1_00_100_000_011_0_x_00;
      patterns[4706] = 33'b1000101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4707] = 33'b1001001101000000_0_1_01_100_000_011_0_x_00;
      patterns[4708] = 33'b1001101101000000_1_1_01_100_000_011_0_x_00;
      patterns[4709] = 33'b1001101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4710] = 33'b1010001101000000_0_1_10_100_000_011_0_x_00;
      patterns[4711] = 33'b1010101101000000_1_1_10_100_000_011_0_x_00;
      patterns[4712] = 33'b1010101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4713] = 33'b1011001101000000_0_1_11_100_000_011_0_x_00;
      patterns[4714] = 33'b1011101101000000_1_1_11_100_000_011_0_x_00;
      patterns[4715] = 33'b1011101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4716] = 33'b0101001101000000_0_1_xx_100_xxx_011_0_1_01;
      patterns[4717] = 33'b0101101101000000_1_1_xx_100_xxx_011_0_1_01;
      patterns[4718] = 33'b0101101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4719] = 33'b0100001101000000_0_0_xx_100_011_xxx_1_x_xx;
      patterns[4720] = 33'b0100101101000000_1_0_xx_100_011_xxx_1_x_xx;
      patterns[4721] = 33'b0100101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4722] = 33'b0000001100001101_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4723] = 33'b0000101100001101_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4724] = 33'b0000101100001101_0_0_00_000_000_000_0_0_00;
      patterns[4725] = 33'b1000001101000001_0_1_00_100_001_011_0_x_00;
      patterns[4726] = 33'b1000101101000001_1_1_00_100_001_011_0_x_00;
      patterns[4727] = 33'b1000101101000001_0_0_00_000_000_000_0_0_00;
      patterns[4728] = 33'b1001001101000001_0_1_01_100_001_011_0_x_00;
      patterns[4729] = 33'b1001101101000001_1_1_01_100_001_011_0_x_00;
      patterns[4730] = 33'b1001101101000001_0_0_00_000_000_000_0_0_00;
      patterns[4731] = 33'b1010001101000001_0_1_10_100_001_011_0_x_00;
      patterns[4732] = 33'b1010101101000001_1_1_10_100_001_011_0_x_00;
      patterns[4733] = 33'b1010101101000001_0_0_00_000_000_000_0_0_00;
      patterns[4734] = 33'b1011001101000001_0_1_11_100_001_011_0_x_00;
      patterns[4735] = 33'b1011101101000001_1_1_11_100_001_011_0_x_00;
      patterns[4736] = 33'b1011101101000001_0_0_00_000_000_000_0_0_00;
      patterns[4737] = 33'b0101001101000000_0_1_xx_100_xxx_011_0_1_01;
      patterns[4738] = 33'b0101101101000000_1_1_xx_100_xxx_011_0_1_01;
      patterns[4739] = 33'b0101101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4740] = 33'b0100001101000000_0_0_xx_100_011_xxx_1_x_xx;
      patterns[4741] = 33'b0100101101000000_1_0_xx_100_011_xxx_1_x_xx;
      patterns[4742] = 33'b0100101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4743] = 33'b0000001100011000_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4744] = 33'b0000101100011000_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4745] = 33'b0000101100011000_0_0_00_000_000_000_0_0_00;
      patterns[4746] = 33'b1000001101000010_0_1_00_100_010_011_0_x_00;
      patterns[4747] = 33'b1000101101000010_1_1_00_100_010_011_0_x_00;
      patterns[4748] = 33'b1000101101000010_0_0_00_000_000_000_0_0_00;
      patterns[4749] = 33'b1001001101000010_0_1_01_100_010_011_0_x_00;
      patterns[4750] = 33'b1001101101000010_1_1_01_100_010_011_0_x_00;
      patterns[4751] = 33'b1001101101000010_0_0_00_000_000_000_0_0_00;
      patterns[4752] = 33'b1010001101000010_0_1_10_100_010_011_0_x_00;
      patterns[4753] = 33'b1010101101000010_1_1_10_100_010_011_0_x_00;
      patterns[4754] = 33'b1010101101000010_0_0_00_000_000_000_0_0_00;
      patterns[4755] = 33'b1011001101000010_0_1_11_100_010_011_0_x_00;
      patterns[4756] = 33'b1011101101000010_1_1_11_100_010_011_0_x_00;
      patterns[4757] = 33'b1011101101000010_0_0_00_000_000_000_0_0_00;
      patterns[4758] = 33'b0101001101000000_0_1_xx_100_xxx_011_0_1_01;
      patterns[4759] = 33'b0101101101000000_1_1_xx_100_xxx_011_0_1_01;
      patterns[4760] = 33'b0101101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4761] = 33'b0100001101000000_0_0_xx_100_011_xxx_1_x_xx;
      patterns[4762] = 33'b0100101101000000_1_0_xx_100_011_xxx_1_x_xx;
      patterns[4763] = 33'b0100101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4764] = 33'b0000001110101111_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4765] = 33'b0000101110101111_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4766] = 33'b0000101110101111_0_0_00_000_000_000_0_0_00;
      patterns[4767] = 33'b1000001101000011_0_1_00_100_011_011_0_x_00;
      patterns[4768] = 33'b1000101101000011_1_1_00_100_011_011_0_x_00;
      patterns[4769] = 33'b1000101101000011_0_0_00_000_000_000_0_0_00;
      patterns[4770] = 33'b1001001101000011_0_1_01_100_011_011_0_x_00;
      patterns[4771] = 33'b1001101101000011_1_1_01_100_011_011_0_x_00;
      patterns[4772] = 33'b1001101101000011_0_0_00_000_000_000_0_0_00;
      patterns[4773] = 33'b1010001101000011_0_1_10_100_011_011_0_x_00;
      patterns[4774] = 33'b1010101101000011_1_1_10_100_011_011_0_x_00;
      patterns[4775] = 33'b1010101101000011_0_0_00_000_000_000_0_0_00;
      patterns[4776] = 33'b1011001101000011_0_1_11_100_011_011_0_x_00;
      patterns[4777] = 33'b1011101101000011_1_1_11_100_011_011_0_x_00;
      patterns[4778] = 33'b1011101101000011_0_0_00_000_000_000_0_0_00;
      patterns[4779] = 33'b0101001101000000_0_1_xx_100_xxx_011_0_1_01;
      patterns[4780] = 33'b0101101101000000_1_1_xx_100_xxx_011_0_1_01;
      patterns[4781] = 33'b0101101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4782] = 33'b0100001101000000_0_0_xx_100_011_xxx_1_x_xx;
      patterns[4783] = 33'b0100101101000000_1_0_xx_100_011_xxx_1_x_xx;
      patterns[4784] = 33'b0100101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4785] = 33'b0000001110000001_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4786] = 33'b0000101110000001_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4787] = 33'b0000101110000001_0_0_00_000_000_000_0_0_00;
      patterns[4788] = 33'b1000001101000100_0_1_00_100_100_011_0_x_00;
      patterns[4789] = 33'b1000101101000100_1_1_00_100_100_011_0_x_00;
      patterns[4790] = 33'b1000101101000100_0_0_00_000_000_000_0_0_00;
      patterns[4791] = 33'b1001001101000100_0_1_01_100_100_011_0_x_00;
      patterns[4792] = 33'b1001101101000100_1_1_01_100_100_011_0_x_00;
      patterns[4793] = 33'b1001101101000100_0_0_00_000_000_000_0_0_00;
      patterns[4794] = 33'b1010001101000100_0_1_10_100_100_011_0_x_00;
      patterns[4795] = 33'b1010101101000100_1_1_10_100_100_011_0_x_00;
      patterns[4796] = 33'b1010101101000100_0_0_00_000_000_000_0_0_00;
      patterns[4797] = 33'b1011001101000100_0_1_11_100_100_011_0_x_00;
      patterns[4798] = 33'b1011101101000100_1_1_11_100_100_011_0_x_00;
      patterns[4799] = 33'b1011101101000100_0_0_00_000_000_000_0_0_00;
      patterns[4800] = 33'b0101001101000000_0_1_xx_100_xxx_011_0_1_01;
      patterns[4801] = 33'b0101101101000000_1_1_xx_100_xxx_011_0_1_01;
      patterns[4802] = 33'b0101101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4803] = 33'b0100001101000000_0_0_xx_100_011_xxx_1_x_xx;
      patterns[4804] = 33'b0100101101000000_1_0_xx_100_011_xxx_1_x_xx;
      patterns[4805] = 33'b0100101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4806] = 33'b0000001101100011_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4807] = 33'b0000101101100011_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4808] = 33'b0000101101100011_0_0_00_000_000_000_0_0_00;
      patterns[4809] = 33'b1000001101000101_0_1_00_100_101_011_0_x_00;
      patterns[4810] = 33'b1000101101000101_1_1_00_100_101_011_0_x_00;
      patterns[4811] = 33'b1000101101000101_0_0_00_000_000_000_0_0_00;
      patterns[4812] = 33'b1001001101000101_0_1_01_100_101_011_0_x_00;
      patterns[4813] = 33'b1001101101000101_1_1_01_100_101_011_0_x_00;
      patterns[4814] = 33'b1001101101000101_0_0_00_000_000_000_0_0_00;
      patterns[4815] = 33'b1010001101000101_0_1_10_100_101_011_0_x_00;
      patterns[4816] = 33'b1010101101000101_1_1_10_100_101_011_0_x_00;
      patterns[4817] = 33'b1010101101000101_0_0_00_000_000_000_0_0_00;
      patterns[4818] = 33'b1011001101000101_0_1_11_100_101_011_0_x_00;
      patterns[4819] = 33'b1011101101000101_1_1_11_100_101_011_0_x_00;
      patterns[4820] = 33'b1011101101000101_0_0_00_000_000_000_0_0_00;
      patterns[4821] = 33'b0101001101000000_0_1_xx_100_xxx_011_0_1_01;
      patterns[4822] = 33'b0101101101000000_1_1_xx_100_xxx_011_0_1_01;
      patterns[4823] = 33'b0101101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4824] = 33'b0100001101000000_0_0_xx_100_011_xxx_1_x_xx;
      patterns[4825] = 33'b0100101101000000_1_0_xx_100_011_xxx_1_x_xx;
      patterns[4826] = 33'b0100101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4827] = 33'b0000001111010110_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4828] = 33'b0000101111010110_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4829] = 33'b0000101111010110_0_0_00_000_000_000_0_0_00;
      patterns[4830] = 33'b1000001101000110_0_1_00_100_110_011_0_x_00;
      patterns[4831] = 33'b1000101101000110_1_1_00_100_110_011_0_x_00;
      patterns[4832] = 33'b1000101101000110_0_0_00_000_000_000_0_0_00;
      patterns[4833] = 33'b1001001101000110_0_1_01_100_110_011_0_x_00;
      patterns[4834] = 33'b1001101101000110_1_1_01_100_110_011_0_x_00;
      patterns[4835] = 33'b1001101101000110_0_0_00_000_000_000_0_0_00;
      patterns[4836] = 33'b1010001101000110_0_1_10_100_110_011_0_x_00;
      patterns[4837] = 33'b1010101101000110_1_1_10_100_110_011_0_x_00;
      patterns[4838] = 33'b1010101101000110_0_0_00_000_000_000_0_0_00;
      patterns[4839] = 33'b1011001101000110_0_1_11_100_110_011_0_x_00;
      patterns[4840] = 33'b1011101101000110_1_1_11_100_110_011_0_x_00;
      patterns[4841] = 33'b1011101101000110_0_0_00_000_000_000_0_0_00;
      patterns[4842] = 33'b0101001101000000_0_1_xx_100_xxx_011_0_1_01;
      patterns[4843] = 33'b0101101101000000_1_1_xx_100_xxx_011_0_1_01;
      patterns[4844] = 33'b0101101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4845] = 33'b0100001101000000_0_0_xx_100_011_xxx_1_x_xx;
      patterns[4846] = 33'b0100101101000000_1_0_xx_100_011_xxx_1_x_xx;
      patterns[4847] = 33'b0100101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4848] = 33'b0000001100010001_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4849] = 33'b0000101100010001_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4850] = 33'b0000101100010001_0_0_00_000_000_000_0_0_00;
      patterns[4851] = 33'b1000001101000111_0_1_00_100_111_011_0_x_00;
      patterns[4852] = 33'b1000101101000111_1_1_00_100_111_011_0_x_00;
      patterns[4853] = 33'b1000101101000111_0_0_00_000_000_000_0_0_00;
      patterns[4854] = 33'b1001001101000111_0_1_01_100_111_011_0_x_00;
      patterns[4855] = 33'b1001101101000111_1_1_01_100_111_011_0_x_00;
      patterns[4856] = 33'b1001101101000111_0_0_00_000_000_000_0_0_00;
      patterns[4857] = 33'b1010001101000111_0_1_10_100_111_011_0_x_00;
      patterns[4858] = 33'b1010101101000111_1_1_10_100_111_011_0_x_00;
      patterns[4859] = 33'b1010101101000111_0_0_00_000_000_000_0_0_00;
      patterns[4860] = 33'b1011001101000111_0_1_11_100_111_011_0_x_00;
      patterns[4861] = 33'b1011101101000111_1_1_11_100_111_011_0_x_00;
      patterns[4862] = 33'b1011101101000111_0_0_00_000_000_000_0_0_00;
      patterns[4863] = 33'b0101001101000000_0_1_xx_100_xxx_011_0_1_01;
      patterns[4864] = 33'b0101101101000000_1_1_xx_100_xxx_011_0_1_01;
      patterns[4865] = 33'b0101101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4866] = 33'b0100001101000000_0_0_xx_100_011_xxx_1_x_xx;
      patterns[4867] = 33'b0100101101000000_1_0_xx_100_011_xxx_1_x_xx;
      patterns[4868] = 33'b0100101101000000_0_0_00_000_000_000_0_0_00;
      patterns[4869] = 33'b0000001100110101_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4870] = 33'b0000101100110101_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4871] = 33'b0000101100110101_0_0_00_000_000_000_0_0_00;
      patterns[4872] = 33'b1000001101010000_0_1_00_101_000_011_0_x_00;
      patterns[4873] = 33'b1000101101010000_1_1_00_101_000_011_0_x_00;
      patterns[4874] = 33'b1000101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4875] = 33'b1001001101010000_0_1_01_101_000_011_0_x_00;
      patterns[4876] = 33'b1001101101010000_1_1_01_101_000_011_0_x_00;
      patterns[4877] = 33'b1001101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4878] = 33'b1010001101010000_0_1_10_101_000_011_0_x_00;
      patterns[4879] = 33'b1010101101010000_1_1_10_101_000_011_0_x_00;
      patterns[4880] = 33'b1010101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4881] = 33'b1011001101010000_0_1_11_101_000_011_0_x_00;
      patterns[4882] = 33'b1011101101010000_1_1_11_101_000_011_0_x_00;
      patterns[4883] = 33'b1011101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4884] = 33'b0101001101010000_0_1_xx_101_xxx_011_0_1_01;
      patterns[4885] = 33'b0101101101010000_1_1_xx_101_xxx_011_0_1_01;
      patterns[4886] = 33'b0101101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4887] = 33'b0100001101010000_0_0_xx_101_011_xxx_1_x_xx;
      patterns[4888] = 33'b0100101101010000_1_0_xx_101_011_xxx_1_x_xx;
      patterns[4889] = 33'b0100101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4890] = 33'b0000001101110001_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4891] = 33'b0000101101110001_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4892] = 33'b0000101101110001_0_0_00_000_000_000_0_0_00;
      patterns[4893] = 33'b1000001101010001_0_1_00_101_001_011_0_x_00;
      patterns[4894] = 33'b1000101101010001_1_1_00_101_001_011_0_x_00;
      patterns[4895] = 33'b1000101101010001_0_0_00_000_000_000_0_0_00;
      patterns[4896] = 33'b1001001101010001_0_1_01_101_001_011_0_x_00;
      patterns[4897] = 33'b1001101101010001_1_1_01_101_001_011_0_x_00;
      patterns[4898] = 33'b1001101101010001_0_0_00_000_000_000_0_0_00;
      patterns[4899] = 33'b1010001101010001_0_1_10_101_001_011_0_x_00;
      patterns[4900] = 33'b1010101101010001_1_1_10_101_001_011_0_x_00;
      patterns[4901] = 33'b1010101101010001_0_0_00_000_000_000_0_0_00;
      patterns[4902] = 33'b1011001101010001_0_1_11_101_001_011_0_x_00;
      patterns[4903] = 33'b1011101101010001_1_1_11_101_001_011_0_x_00;
      patterns[4904] = 33'b1011101101010001_0_0_00_000_000_000_0_0_00;
      patterns[4905] = 33'b0101001101010000_0_1_xx_101_xxx_011_0_1_01;
      patterns[4906] = 33'b0101101101010000_1_1_xx_101_xxx_011_0_1_01;
      patterns[4907] = 33'b0101101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4908] = 33'b0100001101010000_0_0_xx_101_011_xxx_1_x_xx;
      patterns[4909] = 33'b0100101101010000_1_0_xx_101_011_xxx_1_x_xx;
      patterns[4910] = 33'b0100101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4911] = 33'b0000001111100100_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4912] = 33'b0000101111100100_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4913] = 33'b0000101111100100_0_0_00_000_000_000_0_0_00;
      patterns[4914] = 33'b1000001101010010_0_1_00_101_010_011_0_x_00;
      patterns[4915] = 33'b1000101101010010_1_1_00_101_010_011_0_x_00;
      patterns[4916] = 33'b1000101101010010_0_0_00_000_000_000_0_0_00;
      patterns[4917] = 33'b1001001101010010_0_1_01_101_010_011_0_x_00;
      patterns[4918] = 33'b1001101101010010_1_1_01_101_010_011_0_x_00;
      patterns[4919] = 33'b1001101101010010_0_0_00_000_000_000_0_0_00;
      patterns[4920] = 33'b1010001101010010_0_1_10_101_010_011_0_x_00;
      patterns[4921] = 33'b1010101101010010_1_1_10_101_010_011_0_x_00;
      patterns[4922] = 33'b1010101101010010_0_0_00_000_000_000_0_0_00;
      patterns[4923] = 33'b1011001101010010_0_1_11_101_010_011_0_x_00;
      patterns[4924] = 33'b1011101101010010_1_1_11_101_010_011_0_x_00;
      patterns[4925] = 33'b1011101101010010_0_0_00_000_000_000_0_0_00;
      patterns[4926] = 33'b0101001101010000_0_1_xx_101_xxx_011_0_1_01;
      patterns[4927] = 33'b0101101101010000_1_1_xx_101_xxx_011_0_1_01;
      patterns[4928] = 33'b0101101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4929] = 33'b0100001101010000_0_0_xx_101_011_xxx_1_x_xx;
      patterns[4930] = 33'b0100101101010000_1_0_xx_101_011_xxx_1_x_xx;
      patterns[4931] = 33'b0100101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4932] = 33'b0000001100010010_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4933] = 33'b0000101100010010_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4934] = 33'b0000101100010010_0_0_00_000_000_000_0_0_00;
      patterns[4935] = 33'b1000001101010011_0_1_00_101_011_011_0_x_00;
      patterns[4936] = 33'b1000101101010011_1_1_00_101_011_011_0_x_00;
      patterns[4937] = 33'b1000101101010011_0_0_00_000_000_000_0_0_00;
      patterns[4938] = 33'b1001001101010011_0_1_01_101_011_011_0_x_00;
      patterns[4939] = 33'b1001101101010011_1_1_01_101_011_011_0_x_00;
      patterns[4940] = 33'b1001101101010011_0_0_00_000_000_000_0_0_00;
      patterns[4941] = 33'b1010001101010011_0_1_10_101_011_011_0_x_00;
      patterns[4942] = 33'b1010101101010011_1_1_10_101_011_011_0_x_00;
      patterns[4943] = 33'b1010101101010011_0_0_00_000_000_000_0_0_00;
      patterns[4944] = 33'b1011001101010011_0_1_11_101_011_011_0_x_00;
      patterns[4945] = 33'b1011101101010011_1_1_11_101_011_011_0_x_00;
      patterns[4946] = 33'b1011101101010011_0_0_00_000_000_000_0_0_00;
      patterns[4947] = 33'b0101001101010000_0_1_xx_101_xxx_011_0_1_01;
      patterns[4948] = 33'b0101101101010000_1_1_xx_101_xxx_011_0_1_01;
      patterns[4949] = 33'b0101101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4950] = 33'b0100001101010000_0_0_xx_101_011_xxx_1_x_xx;
      patterns[4951] = 33'b0100101101010000_1_0_xx_101_011_xxx_1_x_xx;
      patterns[4952] = 33'b0100101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4953] = 33'b0000001110000001_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4954] = 33'b0000101110000001_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4955] = 33'b0000101110000001_0_0_00_000_000_000_0_0_00;
      patterns[4956] = 33'b1000001101010100_0_1_00_101_100_011_0_x_00;
      patterns[4957] = 33'b1000101101010100_1_1_00_101_100_011_0_x_00;
      patterns[4958] = 33'b1000101101010100_0_0_00_000_000_000_0_0_00;
      patterns[4959] = 33'b1001001101010100_0_1_01_101_100_011_0_x_00;
      patterns[4960] = 33'b1001101101010100_1_1_01_101_100_011_0_x_00;
      patterns[4961] = 33'b1001101101010100_0_0_00_000_000_000_0_0_00;
      patterns[4962] = 33'b1010001101010100_0_1_10_101_100_011_0_x_00;
      patterns[4963] = 33'b1010101101010100_1_1_10_101_100_011_0_x_00;
      patterns[4964] = 33'b1010101101010100_0_0_00_000_000_000_0_0_00;
      patterns[4965] = 33'b1011001101010100_0_1_11_101_100_011_0_x_00;
      patterns[4966] = 33'b1011101101010100_1_1_11_101_100_011_0_x_00;
      patterns[4967] = 33'b1011101101010100_0_0_00_000_000_000_0_0_00;
      patterns[4968] = 33'b0101001101010000_0_1_xx_101_xxx_011_0_1_01;
      patterns[4969] = 33'b0101101101010000_1_1_xx_101_xxx_011_0_1_01;
      patterns[4970] = 33'b0101101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4971] = 33'b0100001101010000_0_0_xx_101_011_xxx_1_x_xx;
      patterns[4972] = 33'b0100101101010000_1_0_xx_101_011_xxx_1_x_xx;
      patterns[4973] = 33'b0100101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4974] = 33'b0000001111000010_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4975] = 33'b0000101111000010_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4976] = 33'b0000101111000010_0_0_00_000_000_000_0_0_00;
      patterns[4977] = 33'b1000001101010101_0_1_00_101_101_011_0_x_00;
      patterns[4978] = 33'b1000101101010101_1_1_00_101_101_011_0_x_00;
      patterns[4979] = 33'b1000101101010101_0_0_00_000_000_000_0_0_00;
      patterns[4980] = 33'b1001001101010101_0_1_01_101_101_011_0_x_00;
      patterns[4981] = 33'b1001101101010101_1_1_01_101_101_011_0_x_00;
      patterns[4982] = 33'b1001101101010101_0_0_00_000_000_000_0_0_00;
      patterns[4983] = 33'b1010001101010101_0_1_10_101_101_011_0_x_00;
      patterns[4984] = 33'b1010101101010101_1_1_10_101_101_011_0_x_00;
      patterns[4985] = 33'b1010101101010101_0_0_00_000_000_000_0_0_00;
      patterns[4986] = 33'b1011001101010101_0_1_11_101_101_011_0_x_00;
      patterns[4987] = 33'b1011101101010101_1_1_11_101_101_011_0_x_00;
      patterns[4988] = 33'b1011101101010101_0_0_00_000_000_000_0_0_00;
      patterns[4989] = 33'b0101001101010000_0_1_xx_101_xxx_011_0_1_01;
      patterns[4990] = 33'b0101101101010000_1_1_xx_101_xxx_011_0_1_01;
      patterns[4991] = 33'b0101101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4992] = 33'b0100001101010000_0_0_xx_101_011_xxx_1_x_xx;
      patterns[4993] = 33'b0100101101010000_1_0_xx_101_011_xxx_1_x_xx;
      patterns[4994] = 33'b0100101101010000_0_0_00_000_000_000_0_0_00;
      patterns[4995] = 33'b0000001111010000_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[4996] = 33'b0000101111010000_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[4997] = 33'b0000101111010000_0_0_00_000_000_000_0_0_00;
      patterns[4998] = 33'b1000001101010110_0_1_00_101_110_011_0_x_00;
      patterns[4999] = 33'b1000101101010110_1_1_00_101_110_011_0_x_00;
      patterns[5000] = 33'b1000101101010110_0_0_00_000_000_000_0_0_00;
      patterns[5001] = 33'b1001001101010110_0_1_01_101_110_011_0_x_00;
      patterns[5002] = 33'b1001101101010110_1_1_01_101_110_011_0_x_00;
      patterns[5003] = 33'b1001101101010110_0_0_00_000_000_000_0_0_00;
      patterns[5004] = 33'b1010001101010110_0_1_10_101_110_011_0_x_00;
      patterns[5005] = 33'b1010101101010110_1_1_10_101_110_011_0_x_00;
      patterns[5006] = 33'b1010101101010110_0_0_00_000_000_000_0_0_00;
      patterns[5007] = 33'b1011001101010110_0_1_11_101_110_011_0_x_00;
      patterns[5008] = 33'b1011101101010110_1_1_11_101_110_011_0_x_00;
      patterns[5009] = 33'b1011101101010110_0_0_00_000_000_000_0_0_00;
      patterns[5010] = 33'b0101001101010000_0_1_xx_101_xxx_011_0_1_01;
      patterns[5011] = 33'b0101101101010000_1_1_xx_101_xxx_011_0_1_01;
      patterns[5012] = 33'b0101101101010000_0_0_00_000_000_000_0_0_00;
      patterns[5013] = 33'b0100001101010000_0_0_xx_101_011_xxx_1_x_xx;
      patterns[5014] = 33'b0100101101010000_1_0_xx_101_011_xxx_1_x_xx;
      patterns[5015] = 33'b0100101101010000_0_0_00_000_000_000_0_0_00;
      patterns[5016] = 33'b0000001100001011_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5017] = 33'b0000101100001011_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5018] = 33'b0000101100001011_0_0_00_000_000_000_0_0_00;
      patterns[5019] = 33'b1000001101010111_0_1_00_101_111_011_0_x_00;
      patterns[5020] = 33'b1000101101010111_1_1_00_101_111_011_0_x_00;
      patterns[5021] = 33'b1000101101010111_0_0_00_000_000_000_0_0_00;
      patterns[5022] = 33'b1001001101010111_0_1_01_101_111_011_0_x_00;
      patterns[5023] = 33'b1001101101010111_1_1_01_101_111_011_0_x_00;
      patterns[5024] = 33'b1001101101010111_0_0_00_000_000_000_0_0_00;
      patterns[5025] = 33'b1010001101010111_0_1_10_101_111_011_0_x_00;
      patterns[5026] = 33'b1010101101010111_1_1_10_101_111_011_0_x_00;
      patterns[5027] = 33'b1010101101010111_0_0_00_000_000_000_0_0_00;
      patterns[5028] = 33'b1011001101010111_0_1_11_101_111_011_0_x_00;
      patterns[5029] = 33'b1011101101010111_1_1_11_101_111_011_0_x_00;
      patterns[5030] = 33'b1011101101010111_0_0_00_000_000_000_0_0_00;
      patterns[5031] = 33'b0101001101010000_0_1_xx_101_xxx_011_0_1_01;
      patterns[5032] = 33'b0101101101010000_1_1_xx_101_xxx_011_0_1_01;
      patterns[5033] = 33'b0101101101010000_0_0_00_000_000_000_0_0_00;
      patterns[5034] = 33'b0100001101010000_0_0_xx_101_011_xxx_1_x_xx;
      patterns[5035] = 33'b0100101101010000_1_0_xx_101_011_xxx_1_x_xx;
      patterns[5036] = 33'b0100101101010000_0_0_00_000_000_000_0_0_00;
      patterns[5037] = 33'b0000001100000101_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5038] = 33'b0000101100000101_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5039] = 33'b0000101100000101_0_0_00_000_000_000_0_0_00;
      patterns[5040] = 33'b1000001101100000_0_1_00_110_000_011_0_x_00;
      patterns[5041] = 33'b1000101101100000_1_1_00_110_000_011_0_x_00;
      patterns[5042] = 33'b1000101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5043] = 33'b1001001101100000_0_1_01_110_000_011_0_x_00;
      patterns[5044] = 33'b1001101101100000_1_1_01_110_000_011_0_x_00;
      patterns[5045] = 33'b1001101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5046] = 33'b1010001101100000_0_1_10_110_000_011_0_x_00;
      patterns[5047] = 33'b1010101101100000_1_1_10_110_000_011_0_x_00;
      patterns[5048] = 33'b1010101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5049] = 33'b1011001101100000_0_1_11_110_000_011_0_x_00;
      patterns[5050] = 33'b1011101101100000_1_1_11_110_000_011_0_x_00;
      patterns[5051] = 33'b1011101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5052] = 33'b0101001101100000_0_1_xx_110_xxx_011_0_1_01;
      patterns[5053] = 33'b0101101101100000_1_1_xx_110_xxx_011_0_1_01;
      patterns[5054] = 33'b0101101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5055] = 33'b0100001101100000_0_0_xx_110_011_xxx_1_x_xx;
      patterns[5056] = 33'b0100101101100000_1_0_xx_110_011_xxx_1_x_xx;
      patterns[5057] = 33'b0100101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5058] = 33'b0000001100011011_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5059] = 33'b0000101100011011_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5060] = 33'b0000101100011011_0_0_00_000_000_000_0_0_00;
      patterns[5061] = 33'b1000001101100001_0_1_00_110_001_011_0_x_00;
      patterns[5062] = 33'b1000101101100001_1_1_00_110_001_011_0_x_00;
      patterns[5063] = 33'b1000101101100001_0_0_00_000_000_000_0_0_00;
      patterns[5064] = 33'b1001001101100001_0_1_01_110_001_011_0_x_00;
      patterns[5065] = 33'b1001101101100001_1_1_01_110_001_011_0_x_00;
      patterns[5066] = 33'b1001101101100001_0_0_00_000_000_000_0_0_00;
      patterns[5067] = 33'b1010001101100001_0_1_10_110_001_011_0_x_00;
      patterns[5068] = 33'b1010101101100001_1_1_10_110_001_011_0_x_00;
      patterns[5069] = 33'b1010101101100001_0_0_00_000_000_000_0_0_00;
      patterns[5070] = 33'b1011001101100001_0_1_11_110_001_011_0_x_00;
      patterns[5071] = 33'b1011101101100001_1_1_11_110_001_011_0_x_00;
      patterns[5072] = 33'b1011101101100001_0_0_00_000_000_000_0_0_00;
      patterns[5073] = 33'b0101001101100000_0_1_xx_110_xxx_011_0_1_01;
      patterns[5074] = 33'b0101101101100000_1_1_xx_110_xxx_011_0_1_01;
      patterns[5075] = 33'b0101101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5076] = 33'b0100001101100000_0_0_xx_110_011_xxx_1_x_xx;
      patterns[5077] = 33'b0100101101100000_1_0_xx_110_011_xxx_1_x_xx;
      patterns[5078] = 33'b0100101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5079] = 33'b0000001110000010_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5080] = 33'b0000101110000010_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5081] = 33'b0000101110000010_0_0_00_000_000_000_0_0_00;
      patterns[5082] = 33'b1000001101100010_0_1_00_110_010_011_0_x_00;
      patterns[5083] = 33'b1000101101100010_1_1_00_110_010_011_0_x_00;
      patterns[5084] = 33'b1000101101100010_0_0_00_000_000_000_0_0_00;
      patterns[5085] = 33'b1001001101100010_0_1_01_110_010_011_0_x_00;
      patterns[5086] = 33'b1001101101100010_1_1_01_110_010_011_0_x_00;
      patterns[5087] = 33'b1001101101100010_0_0_00_000_000_000_0_0_00;
      patterns[5088] = 33'b1010001101100010_0_1_10_110_010_011_0_x_00;
      patterns[5089] = 33'b1010101101100010_1_1_10_110_010_011_0_x_00;
      patterns[5090] = 33'b1010101101100010_0_0_00_000_000_000_0_0_00;
      patterns[5091] = 33'b1011001101100010_0_1_11_110_010_011_0_x_00;
      patterns[5092] = 33'b1011101101100010_1_1_11_110_010_011_0_x_00;
      patterns[5093] = 33'b1011101101100010_0_0_00_000_000_000_0_0_00;
      patterns[5094] = 33'b0101001101100000_0_1_xx_110_xxx_011_0_1_01;
      patterns[5095] = 33'b0101101101100000_1_1_xx_110_xxx_011_0_1_01;
      patterns[5096] = 33'b0101101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5097] = 33'b0100001101100000_0_0_xx_110_011_xxx_1_x_xx;
      patterns[5098] = 33'b0100101101100000_1_0_xx_110_011_xxx_1_x_xx;
      patterns[5099] = 33'b0100101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5100] = 33'b0000001110010110_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5101] = 33'b0000101110010110_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5102] = 33'b0000101110010110_0_0_00_000_000_000_0_0_00;
      patterns[5103] = 33'b1000001101100011_0_1_00_110_011_011_0_x_00;
      patterns[5104] = 33'b1000101101100011_1_1_00_110_011_011_0_x_00;
      patterns[5105] = 33'b1000101101100011_0_0_00_000_000_000_0_0_00;
      patterns[5106] = 33'b1001001101100011_0_1_01_110_011_011_0_x_00;
      patterns[5107] = 33'b1001101101100011_1_1_01_110_011_011_0_x_00;
      patterns[5108] = 33'b1001101101100011_0_0_00_000_000_000_0_0_00;
      patterns[5109] = 33'b1010001101100011_0_1_10_110_011_011_0_x_00;
      patterns[5110] = 33'b1010101101100011_1_1_10_110_011_011_0_x_00;
      patterns[5111] = 33'b1010101101100011_0_0_00_000_000_000_0_0_00;
      patterns[5112] = 33'b1011001101100011_0_1_11_110_011_011_0_x_00;
      patterns[5113] = 33'b1011101101100011_1_1_11_110_011_011_0_x_00;
      patterns[5114] = 33'b1011101101100011_0_0_00_000_000_000_0_0_00;
      patterns[5115] = 33'b0101001101100000_0_1_xx_110_xxx_011_0_1_01;
      patterns[5116] = 33'b0101101101100000_1_1_xx_110_xxx_011_0_1_01;
      patterns[5117] = 33'b0101101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5118] = 33'b0100001101100000_0_0_xx_110_011_xxx_1_x_xx;
      patterns[5119] = 33'b0100101101100000_1_0_xx_110_011_xxx_1_x_xx;
      patterns[5120] = 33'b0100101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5121] = 33'b0000001101001111_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5122] = 33'b0000101101001111_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5123] = 33'b0000101101001111_0_0_00_000_000_000_0_0_00;
      patterns[5124] = 33'b1000001101100100_0_1_00_110_100_011_0_x_00;
      patterns[5125] = 33'b1000101101100100_1_1_00_110_100_011_0_x_00;
      patterns[5126] = 33'b1000101101100100_0_0_00_000_000_000_0_0_00;
      patterns[5127] = 33'b1001001101100100_0_1_01_110_100_011_0_x_00;
      patterns[5128] = 33'b1001101101100100_1_1_01_110_100_011_0_x_00;
      patterns[5129] = 33'b1001101101100100_0_0_00_000_000_000_0_0_00;
      patterns[5130] = 33'b1010001101100100_0_1_10_110_100_011_0_x_00;
      patterns[5131] = 33'b1010101101100100_1_1_10_110_100_011_0_x_00;
      patterns[5132] = 33'b1010101101100100_0_0_00_000_000_000_0_0_00;
      patterns[5133] = 33'b1011001101100100_0_1_11_110_100_011_0_x_00;
      patterns[5134] = 33'b1011101101100100_1_1_11_110_100_011_0_x_00;
      patterns[5135] = 33'b1011101101100100_0_0_00_000_000_000_0_0_00;
      patterns[5136] = 33'b0101001101100000_0_1_xx_110_xxx_011_0_1_01;
      patterns[5137] = 33'b0101101101100000_1_1_xx_110_xxx_011_0_1_01;
      patterns[5138] = 33'b0101101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5139] = 33'b0100001101100000_0_0_xx_110_011_xxx_1_x_xx;
      patterns[5140] = 33'b0100101101100000_1_0_xx_110_011_xxx_1_x_xx;
      patterns[5141] = 33'b0100101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5142] = 33'b0000001111110111_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5143] = 33'b0000101111110111_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5144] = 33'b0000101111110111_0_0_00_000_000_000_0_0_00;
      patterns[5145] = 33'b1000001101100101_0_1_00_110_101_011_0_x_00;
      patterns[5146] = 33'b1000101101100101_1_1_00_110_101_011_0_x_00;
      patterns[5147] = 33'b1000101101100101_0_0_00_000_000_000_0_0_00;
      patterns[5148] = 33'b1001001101100101_0_1_01_110_101_011_0_x_00;
      patterns[5149] = 33'b1001101101100101_1_1_01_110_101_011_0_x_00;
      patterns[5150] = 33'b1001101101100101_0_0_00_000_000_000_0_0_00;
      patterns[5151] = 33'b1010001101100101_0_1_10_110_101_011_0_x_00;
      patterns[5152] = 33'b1010101101100101_1_1_10_110_101_011_0_x_00;
      patterns[5153] = 33'b1010101101100101_0_0_00_000_000_000_0_0_00;
      patterns[5154] = 33'b1011001101100101_0_1_11_110_101_011_0_x_00;
      patterns[5155] = 33'b1011101101100101_1_1_11_110_101_011_0_x_00;
      patterns[5156] = 33'b1011101101100101_0_0_00_000_000_000_0_0_00;
      patterns[5157] = 33'b0101001101100000_0_1_xx_110_xxx_011_0_1_01;
      patterns[5158] = 33'b0101101101100000_1_1_xx_110_xxx_011_0_1_01;
      patterns[5159] = 33'b0101101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5160] = 33'b0100001101100000_0_0_xx_110_011_xxx_1_x_xx;
      patterns[5161] = 33'b0100101101100000_1_0_xx_110_011_xxx_1_x_xx;
      patterns[5162] = 33'b0100101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5163] = 33'b0000001101000010_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5164] = 33'b0000101101000010_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5165] = 33'b0000101101000010_0_0_00_000_000_000_0_0_00;
      patterns[5166] = 33'b1000001101100110_0_1_00_110_110_011_0_x_00;
      patterns[5167] = 33'b1000101101100110_1_1_00_110_110_011_0_x_00;
      patterns[5168] = 33'b1000101101100110_0_0_00_000_000_000_0_0_00;
      patterns[5169] = 33'b1001001101100110_0_1_01_110_110_011_0_x_00;
      patterns[5170] = 33'b1001101101100110_1_1_01_110_110_011_0_x_00;
      patterns[5171] = 33'b1001101101100110_0_0_00_000_000_000_0_0_00;
      patterns[5172] = 33'b1010001101100110_0_1_10_110_110_011_0_x_00;
      patterns[5173] = 33'b1010101101100110_1_1_10_110_110_011_0_x_00;
      patterns[5174] = 33'b1010101101100110_0_0_00_000_000_000_0_0_00;
      patterns[5175] = 33'b1011001101100110_0_1_11_110_110_011_0_x_00;
      patterns[5176] = 33'b1011101101100110_1_1_11_110_110_011_0_x_00;
      patterns[5177] = 33'b1011101101100110_0_0_00_000_000_000_0_0_00;
      patterns[5178] = 33'b0101001101100000_0_1_xx_110_xxx_011_0_1_01;
      patterns[5179] = 33'b0101101101100000_1_1_xx_110_xxx_011_0_1_01;
      patterns[5180] = 33'b0101101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5181] = 33'b0100001101100000_0_0_xx_110_011_xxx_1_x_xx;
      patterns[5182] = 33'b0100101101100000_1_0_xx_110_011_xxx_1_x_xx;
      patterns[5183] = 33'b0100101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5184] = 33'b0000001111001111_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5185] = 33'b0000101111001111_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5186] = 33'b0000101111001111_0_0_00_000_000_000_0_0_00;
      patterns[5187] = 33'b1000001101100111_0_1_00_110_111_011_0_x_00;
      patterns[5188] = 33'b1000101101100111_1_1_00_110_111_011_0_x_00;
      patterns[5189] = 33'b1000101101100111_0_0_00_000_000_000_0_0_00;
      patterns[5190] = 33'b1001001101100111_0_1_01_110_111_011_0_x_00;
      patterns[5191] = 33'b1001101101100111_1_1_01_110_111_011_0_x_00;
      patterns[5192] = 33'b1001101101100111_0_0_00_000_000_000_0_0_00;
      patterns[5193] = 33'b1010001101100111_0_1_10_110_111_011_0_x_00;
      patterns[5194] = 33'b1010101101100111_1_1_10_110_111_011_0_x_00;
      patterns[5195] = 33'b1010101101100111_0_0_00_000_000_000_0_0_00;
      patterns[5196] = 33'b1011001101100111_0_1_11_110_111_011_0_x_00;
      patterns[5197] = 33'b1011101101100111_1_1_11_110_111_011_0_x_00;
      patterns[5198] = 33'b1011101101100111_0_0_00_000_000_000_0_0_00;
      patterns[5199] = 33'b0101001101100000_0_1_xx_110_xxx_011_0_1_01;
      patterns[5200] = 33'b0101101101100000_1_1_xx_110_xxx_011_0_1_01;
      patterns[5201] = 33'b0101101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5202] = 33'b0100001101100000_0_0_xx_110_011_xxx_1_x_xx;
      patterns[5203] = 33'b0100101101100000_1_0_xx_110_011_xxx_1_x_xx;
      patterns[5204] = 33'b0100101101100000_0_0_00_000_000_000_0_0_00;
      patterns[5205] = 33'b0000001110001111_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5206] = 33'b0000101110001111_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5207] = 33'b0000101110001111_0_0_00_000_000_000_0_0_00;
      patterns[5208] = 33'b1000001101110000_0_1_00_111_000_011_0_x_00;
      patterns[5209] = 33'b1000101101110000_1_1_00_111_000_011_0_x_00;
      patterns[5210] = 33'b1000101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5211] = 33'b1001001101110000_0_1_01_111_000_011_0_x_00;
      patterns[5212] = 33'b1001101101110000_1_1_01_111_000_011_0_x_00;
      patterns[5213] = 33'b1001101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5214] = 33'b1010001101110000_0_1_10_111_000_011_0_x_00;
      patterns[5215] = 33'b1010101101110000_1_1_10_111_000_011_0_x_00;
      patterns[5216] = 33'b1010101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5217] = 33'b1011001101110000_0_1_11_111_000_011_0_x_00;
      patterns[5218] = 33'b1011101101110000_1_1_11_111_000_011_0_x_00;
      patterns[5219] = 33'b1011101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5220] = 33'b0101001101110000_0_1_xx_111_xxx_011_0_1_01;
      patterns[5221] = 33'b0101101101110000_1_1_xx_111_xxx_011_0_1_01;
      patterns[5222] = 33'b0101101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5223] = 33'b0100001101110000_0_0_xx_111_011_xxx_1_x_xx;
      patterns[5224] = 33'b0100101101110000_1_0_xx_111_011_xxx_1_x_xx;
      patterns[5225] = 33'b0100101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5226] = 33'b0000001101111111_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5227] = 33'b0000101101111111_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5228] = 33'b0000101101111111_0_0_00_000_000_000_0_0_00;
      patterns[5229] = 33'b1000001101110001_0_1_00_111_001_011_0_x_00;
      patterns[5230] = 33'b1000101101110001_1_1_00_111_001_011_0_x_00;
      patterns[5231] = 33'b1000101101110001_0_0_00_000_000_000_0_0_00;
      patterns[5232] = 33'b1001001101110001_0_1_01_111_001_011_0_x_00;
      patterns[5233] = 33'b1001101101110001_1_1_01_111_001_011_0_x_00;
      patterns[5234] = 33'b1001101101110001_0_0_00_000_000_000_0_0_00;
      patterns[5235] = 33'b1010001101110001_0_1_10_111_001_011_0_x_00;
      patterns[5236] = 33'b1010101101110001_1_1_10_111_001_011_0_x_00;
      patterns[5237] = 33'b1010101101110001_0_0_00_000_000_000_0_0_00;
      patterns[5238] = 33'b1011001101110001_0_1_11_111_001_011_0_x_00;
      patterns[5239] = 33'b1011101101110001_1_1_11_111_001_011_0_x_00;
      patterns[5240] = 33'b1011101101110001_0_0_00_000_000_000_0_0_00;
      patterns[5241] = 33'b0101001101110000_0_1_xx_111_xxx_011_0_1_01;
      patterns[5242] = 33'b0101101101110000_1_1_xx_111_xxx_011_0_1_01;
      patterns[5243] = 33'b0101101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5244] = 33'b0100001101110000_0_0_xx_111_011_xxx_1_x_xx;
      patterns[5245] = 33'b0100101101110000_1_0_xx_111_011_xxx_1_x_xx;
      patterns[5246] = 33'b0100101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5247] = 33'b0000001111001110_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5248] = 33'b0000101111001110_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5249] = 33'b0000101111001110_0_0_00_000_000_000_0_0_00;
      patterns[5250] = 33'b1000001101110010_0_1_00_111_010_011_0_x_00;
      patterns[5251] = 33'b1000101101110010_1_1_00_111_010_011_0_x_00;
      patterns[5252] = 33'b1000101101110010_0_0_00_000_000_000_0_0_00;
      patterns[5253] = 33'b1001001101110010_0_1_01_111_010_011_0_x_00;
      patterns[5254] = 33'b1001101101110010_1_1_01_111_010_011_0_x_00;
      patterns[5255] = 33'b1001101101110010_0_0_00_000_000_000_0_0_00;
      patterns[5256] = 33'b1010001101110010_0_1_10_111_010_011_0_x_00;
      patterns[5257] = 33'b1010101101110010_1_1_10_111_010_011_0_x_00;
      patterns[5258] = 33'b1010101101110010_0_0_00_000_000_000_0_0_00;
      patterns[5259] = 33'b1011001101110010_0_1_11_111_010_011_0_x_00;
      patterns[5260] = 33'b1011101101110010_1_1_11_111_010_011_0_x_00;
      patterns[5261] = 33'b1011101101110010_0_0_00_000_000_000_0_0_00;
      patterns[5262] = 33'b0101001101110000_0_1_xx_111_xxx_011_0_1_01;
      patterns[5263] = 33'b0101101101110000_1_1_xx_111_xxx_011_0_1_01;
      patterns[5264] = 33'b0101101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5265] = 33'b0100001101110000_0_0_xx_111_011_xxx_1_x_xx;
      patterns[5266] = 33'b0100101101110000_1_0_xx_111_011_xxx_1_x_xx;
      patterns[5267] = 33'b0100101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5268] = 33'b0000001101010111_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5269] = 33'b0000101101010111_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5270] = 33'b0000101101010111_0_0_00_000_000_000_0_0_00;
      patterns[5271] = 33'b1000001101110011_0_1_00_111_011_011_0_x_00;
      patterns[5272] = 33'b1000101101110011_1_1_00_111_011_011_0_x_00;
      patterns[5273] = 33'b1000101101110011_0_0_00_000_000_000_0_0_00;
      patterns[5274] = 33'b1001001101110011_0_1_01_111_011_011_0_x_00;
      patterns[5275] = 33'b1001101101110011_1_1_01_111_011_011_0_x_00;
      patterns[5276] = 33'b1001101101110011_0_0_00_000_000_000_0_0_00;
      patterns[5277] = 33'b1010001101110011_0_1_10_111_011_011_0_x_00;
      patterns[5278] = 33'b1010101101110011_1_1_10_111_011_011_0_x_00;
      patterns[5279] = 33'b1010101101110011_0_0_00_000_000_000_0_0_00;
      patterns[5280] = 33'b1011001101110011_0_1_11_111_011_011_0_x_00;
      patterns[5281] = 33'b1011101101110011_1_1_11_111_011_011_0_x_00;
      patterns[5282] = 33'b1011101101110011_0_0_00_000_000_000_0_0_00;
      patterns[5283] = 33'b0101001101110000_0_1_xx_111_xxx_011_0_1_01;
      patterns[5284] = 33'b0101101101110000_1_1_xx_111_xxx_011_0_1_01;
      patterns[5285] = 33'b0101101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5286] = 33'b0100001101110000_0_0_xx_111_011_xxx_1_x_xx;
      patterns[5287] = 33'b0100101101110000_1_0_xx_111_011_xxx_1_x_xx;
      patterns[5288] = 33'b0100101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5289] = 33'b0000001110000100_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5290] = 33'b0000101110000100_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5291] = 33'b0000101110000100_0_0_00_000_000_000_0_0_00;
      patterns[5292] = 33'b1000001101110100_0_1_00_111_100_011_0_x_00;
      patterns[5293] = 33'b1000101101110100_1_1_00_111_100_011_0_x_00;
      patterns[5294] = 33'b1000101101110100_0_0_00_000_000_000_0_0_00;
      patterns[5295] = 33'b1001001101110100_0_1_01_111_100_011_0_x_00;
      patterns[5296] = 33'b1001101101110100_1_1_01_111_100_011_0_x_00;
      patterns[5297] = 33'b1001101101110100_0_0_00_000_000_000_0_0_00;
      patterns[5298] = 33'b1010001101110100_0_1_10_111_100_011_0_x_00;
      patterns[5299] = 33'b1010101101110100_1_1_10_111_100_011_0_x_00;
      patterns[5300] = 33'b1010101101110100_0_0_00_000_000_000_0_0_00;
      patterns[5301] = 33'b1011001101110100_0_1_11_111_100_011_0_x_00;
      patterns[5302] = 33'b1011101101110100_1_1_11_111_100_011_0_x_00;
      patterns[5303] = 33'b1011101101110100_0_0_00_000_000_000_0_0_00;
      patterns[5304] = 33'b0101001101110000_0_1_xx_111_xxx_011_0_1_01;
      patterns[5305] = 33'b0101101101110000_1_1_xx_111_xxx_011_0_1_01;
      patterns[5306] = 33'b0101101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5307] = 33'b0100001101110000_0_0_xx_111_011_xxx_1_x_xx;
      patterns[5308] = 33'b0100101101110000_1_0_xx_111_011_xxx_1_x_xx;
      patterns[5309] = 33'b0100101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5310] = 33'b0000001100100110_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5311] = 33'b0000101100100110_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5312] = 33'b0000101100100110_0_0_00_000_000_000_0_0_00;
      patterns[5313] = 33'b1000001101110101_0_1_00_111_101_011_0_x_00;
      patterns[5314] = 33'b1000101101110101_1_1_00_111_101_011_0_x_00;
      patterns[5315] = 33'b1000101101110101_0_0_00_000_000_000_0_0_00;
      patterns[5316] = 33'b1001001101110101_0_1_01_111_101_011_0_x_00;
      patterns[5317] = 33'b1001101101110101_1_1_01_111_101_011_0_x_00;
      patterns[5318] = 33'b1001101101110101_0_0_00_000_000_000_0_0_00;
      patterns[5319] = 33'b1010001101110101_0_1_10_111_101_011_0_x_00;
      patterns[5320] = 33'b1010101101110101_1_1_10_111_101_011_0_x_00;
      patterns[5321] = 33'b1010101101110101_0_0_00_000_000_000_0_0_00;
      patterns[5322] = 33'b1011001101110101_0_1_11_111_101_011_0_x_00;
      patterns[5323] = 33'b1011101101110101_1_1_11_111_101_011_0_x_00;
      patterns[5324] = 33'b1011101101110101_0_0_00_000_000_000_0_0_00;
      patterns[5325] = 33'b0101001101110000_0_1_xx_111_xxx_011_0_1_01;
      patterns[5326] = 33'b0101101101110000_1_1_xx_111_xxx_011_0_1_01;
      patterns[5327] = 33'b0101101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5328] = 33'b0100001101110000_0_0_xx_111_011_xxx_1_x_xx;
      patterns[5329] = 33'b0100101101110000_1_0_xx_111_011_xxx_1_x_xx;
      patterns[5330] = 33'b0100101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5331] = 33'b0000001101111101_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5332] = 33'b0000101101111101_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5333] = 33'b0000101101111101_0_0_00_000_000_000_0_0_00;
      patterns[5334] = 33'b1000001101110110_0_1_00_111_110_011_0_x_00;
      patterns[5335] = 33'b1000101101110110_1_1_00_111_110_011_0_x_00;
      patterns[5336] = 33'b1000101101110110_0_0_00_000_000_000_0_0_00;
      patterns[5337] = 33'b1001001101110110_0_1_01_111_110_011_0_x_00;
      patterns[5338] = 33'b1001101101110110_1_1_01_111_110_011_0_x_00;
      patterns[5339] = 33'b1001101101110110_0_0_00_000_000_000_0_0_00;
      patterns[5340] = 33'b1010001101110110_0_1_10_111_110_011_0_x_00;
      patterns[5341] = 33'b1010101101110110_1_1_10_111_110_011_0_x_00;
      patterns[5342] = 33'b1010101101110110_0_0_00_000_000_000_0_0_00;
      patterns[5343] = 33'b1011001101110110_0_1_11_111_110_011_0_x_00;
      patterns[5344] = 33'b1011101101110110_1_1_11_111_110_011_0_x_00;
      patterns[5345] = 33'b1011101101110110_0_0_00_000_000_000_0_0_00;
      patterns[5346] = 33'b0101001101110000_0_1_xx_111_xxx_011_0_1_01;
      patterns[5347] = 33'b0101101101110000_1_1_xx_111_xxx_011_0_1_01;
      patterns[5348] = 33'b0101101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5349] = 33'b0100001101110000_0_0_xx_111_011_xxx_1_x_xx;
      patterns[5350] = 33'b0100101101110000_1_0_xx_111_011_xxx_1_x_xx;
      patterns[5351] = 33'b0100101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5352] = 33'b0000001100011101_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5353] = 33'b0000101100011101_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5354] = 33'b0000101100011101_0_0_00_000_000_000_0_0_00;
      patterns[5355] = 33'b1000001101110111_0_1_00_111_111_011_0_x_00;
      patterns[5356] = 33'b1000101101110111_1_1_00_111_111_011_0_x_00;
      patterns[5357] = 33'b1000101101110111_0_0_00_000_000_000_0_0_00;
      patterns[5358] = 33'b1001001101110111_0_1_01_111_111_011_0_x_00;
      patterns[5359] = 33'b1001101101110111_1_1_01_111_111_011_0_x_00;
      patterns[5360] = 33'b1001101101110111_0_0_00_000_000_000_0_0_00;
      patterns[5361] = 33'b1010001101110111_0_1_10_111_111_011_0_x_00;
      patterns[5362] = 33'b1010101101110111_1_1_10_111_111_011_0_x_00;
      patterns[5363] = 33'b1010101101110111_0_0_00_000_000_000_0_0_00;
      patterns[5364] = 33'b1011001101110111_0_1_11_111_111_011_0_x_00;
      patterns[5365] = 33'b1011101101110111_1_1_11_111_111_011_0_x_00;
      patterns[5366] = 33'b1011101101110111_0_0_00_000_000_000_0_0_00;
      patterns[5367] = 33'b0101001101110000_0_1_xx_111_xxx_011_0_1_01;
      patterns[5368] = 33'b0101101101110000_1_1_xx_111_xxx_011_0_1_01;
      patterns[5369] = 33'b0101101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5370] = 33'b0100001101110000_0_0_xx_111_011_xxx_1_x_xx;
      patterns[5371] = 33'b0100101101110000_1_0_xx_111_011_xxx_1_x_xx;
      patterns[5372] = 33'b0100101101110000_0_0_00_000_000_000_0_0_00;
      patterns[5373] = 33'b0000001101010110_0_1_xx_xxx_xxx_011_0_x_10;
      patterns[5374] = 33'b0000101101010110_1_1_xx_xxx_xxx_011_0_x_10;
      patterns[5375] = 33'b0000101101010110_0_0_00_000_000_000_0_0_00;
      patterns[5376] = 33'b1000010000000000_0_1_00_000_000_100_0_x_00;
      patterns[5377] = 33'b1000110000000000_1_1_00_000_000_100_0_x_00;
      patterns[5378] = 33'b1000110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5379] = 33'b1001010000000000_0_1_01_000_000_100_0_x_00;
      patterns[5380] = 33'b1001110000000000_1_1_01_000_000_100_0_x_00;
      patterns[5381] = 33'b1001110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5382] = 33'b1010010000000000_0_1_10_000_000_100_0_x_00;
      patterns[5383] = 33'b1010110000000000_1_1_10_000_000_100_0_x_00;
      patterns[5384] = 33'b1010110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5385] = 33'b1011010000000000_0_1_11_000_000_100_0_x_00;
      patterns[5386] = 33'b1011110000000000_1_1_11_000_000_100_0_x_00;
      patterns[5387] = 33'b1011110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5388] = 33'b0101010000000000_0_1_xx_000_xxx_100_0_1_01;
      patterns[5389] = 33'b0101110000000000_1_1_xx_000_xxx_100_0_1_01;
      patterns[5390] = 33'b0101110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5391] = 33'b0100010000000000_0_0_xx_000_100_xxx_1_x_xx;
      patterns[5392] = 33'b0100110000000000_1_0_xx_000_100_xxx_1_x_xx;
      patterns[5393] = 33'b0100110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5394] = 33'b0000010000000111_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5395] = 33'b0000110000000111_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5396] = 33'b0000110000000111_0_0_00_000_000_000_0_0_00;
      patterns[5397] = 33'b1000010000000001_0_1_00_000_001_100_0_x_00;
      patterns[5398] = 33'b1000110000000001_1_1_00_000_001_100_0_x_00;
      patterns[5399] = 33'b1000110000000001_0_0_00_000_000_000_0_0_00;
      patterns[5400] = 33'b1001010000000001_0_1_01_000_001_100_0_x_00;
      patterns[5401] = 33'b1001110000000001_1_1_01_000_001_100_0_x_00;
      patterns[5402] = 33'b1001110000000001_0_0_00_000_000_000_0_0_00;
      patterns[5403] = 33'b1010010000000001_0_1_10_000_001_100_0_x_00;
      patterns[5404] = 33'b1010110000000001_1_1_10_000_001_100_0_x_00;
      patterns[5405] = 33'b1010110000000001_0_0_00_000_000_000_0_0_00;
      patterns[5406] = 33'b1011010000000001_0_1_11_000_001_100_0_x_00;
      patterns[5407] = 33'b1011110000000001_1_1_11_000_001_100_0_x_00;
      patterns[5408] = 33'b1011110000000001_0_0_00_000_000_000_0_0_00;
      patterns[5409] = 33'b0101010000000000_0_1_xx_000_xxx_100_0_1_01;
      patterns[5410] = 33'b0101110000000000_1_1_xx_000_xxx_100_0_1_01;
      patterns[5411] = 33'b0101110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5412] = 33'b0100010000000000_0_0_xx_000_100_xxx_1_x_xx;
      patterns[5413] = 33'b0100110000000000_1_0_xx_000_100_xxx_1_x_xx;
      patterns[5414] = 33'b0100110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5415] = 33'b0000010000101100_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5416] = 33'b0000110000101100_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5417] = 33'b0000110000101100_0_0_00_000_000_000_0_0_00;
      patterns[5418] = 33'b1000010000000010_0_1_00_000_010_100_0_x_00;
      patterns[5419] = 33'b1000110000000010_1_1_00_000_010_100_0_x_00;
      patterns[5420] = 33'b1000110000000010_0_0_00_000_000_000_0_0_00;
      patterns[5421] = 33'b1001010000000010_0_1_01_000_010_100_0_x_00;
      patterns[5422] = 33'b1001110000000010_1_1_01_000_010_100_0_x_00;
      patterns[5423] = 33'b1001110000000010_0_0_00_000_000_000_0_0_00;
      patterns[5424] = 33'b1010010000000010_0_1_10_000_010_100_0_x_00;
      patterns[5425] = 33'b1010110000000010_1_1_10_000_010_100_0_x_00;
      patterns[5426] = 33'b1010110000000010_0_0_00_000_000_000_0_0_00;
      patterns[5427] = 33'b1011010000000010_0_1_11_000_010_100_0_x_00;
      patterns[5428] = 33'b1011110000000010_1_1_11_000_010_100_0_x_00;
      patterns[5429] = 33'b1011110000000010_0_0_00_000_000_000_0_0_00;
      patterns[5430] = 33'b0101010000000000_0_1_xx_000_xxx_100_0_1_01;
      patterns[5431] = 33'b0101110000000000_1_1_xx_000_xxx_100_0_1_01;
      patterns[5432] = 33'b0101110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5433] = 33'b0100010000000000_0_0_xx_000_100_xxx_1_x_xx;
      patterns[5434] = 33'b0100110000000000_1_0_xx_000_100_xxx_1_x_xx;
      patterns[5435] = 33'b0100110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5436] = 33'b0000010000101000_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5437] = 33'b0000110000101000_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5438] = 33'b0000110000101000_0_0_00_000_000_000_0_0_00;
      patterns[5439] = 33'b1000010000000011_0_1_00_000_011_100_0_x_00;
      patterns[5440] = 33'b1000110000000011_1_1_00_000_011_100_0_x_00;
      patterns[5441] = 33'b1000110000000011_0_0_00_000_000_000_0_0_00;
      patterns[5442] = 33'b1001010000000011_0_1_01_000_011_100_0_x_00;
      patterns[5443] = 33'b1001110000000011_1_1_01_000_011_100_0_x_00;
      patterns[5444] = 33'b1001110000000011_0_0_00_000_000_000_0_0_00;
      patterns[5445] = 33'b1010010000000011_0_1_10_000_011_100_0_x_00;
      patterns[5446] = 33'b1010110000000011_1_1_10_000_011_100_0_x_00;
      patterns[5447] = 33'b1010110000000011_0_0_00_000_000_000_0_0_00;
      patterns[5448] = 33'b1011010000000011_0_1_11_000_011_100_0_x_00;
      patterns[5449] = 33'b1011110000000011_1_1_11_000_011_100_0_x_00;
      patterns[5450] = 33'b1011110000000011_0_0_00_000_000_000_0_0_00;
      patterns[5451] = 33'b0101010000000000_0_1_xx_000_xxx_100_0_1_01;
      patterns[5452] = 33'b0101110000000000_1_1_xx_000_xxx_100_0_1_01;
      patterns[5453] = 33'b0101110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5454] = 33'b0100010000000000_0_0_xx_000_100_xxx_1_x_xx;
      patterns[5455] = 33'b0100110000000000_1_0_xx_000_100_xxx_1_x_xx;
      patterns[5456] = 33'b0100110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5457] = 33'b0000010001111110_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5458] = 33'b0000110001111110_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5459] = 33'b0000110001111110_0_0_00_000_000_000_0_0_00;
      patterns[5460] = 33'b1000010000000100_0_1_00_000_100_100_0_x_00;
      patterns[5461] = 33'b1000110000000100_1_1_00_000_100_100_0_x_00;
      patterns[5462] = 33'b1000110000000100_0_0_00_000_000_000_0_0_00;
      patterns[5463] = 33'b1001010000000100_0_1_01_000_100_100_0_x_00;
      patterns[5464] = 33'b1001110000000100_1_1_01_000_100_100_0_x_00;
      patterns[5465] = 33'b1001110000000100_0_0_00_000_000_000_0_0_00;
      patterns[5466] = 33'b1010010000000100_0_1_10_000_100_100_0_x_00;
      patterns[5467] = 33'b1010110000000100_1_1_10_000_100_100_0_x_00;
      patterns[5468] = 33'b1010110000000100_0_0_00_000_000_000_0_0_00;
      patterns[5469] = 33'b1011010000000100_0_1_11_000_100_100_0_x_00;
      patterns[5470] = 33'b1011110000000100_1_1_11_000_100_100_0_x_00;
      patterns[5471] = 33'b1011110000000100_0_0_00_000_000_000_0_0_00;
      patterns[5472] = 33'b0101010000000000_0_1_xx_000_xxx_100_0_1_01;
      patterns[5473] = 33'b0101110000000000_1_1_xx_000_xxx_100_0_1_01;
      patterns[5474] = 33'b0101110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5475] = 33'b0100010000000000_0_0_xx_000_100_xxx_1_x_xx;
      patterns[5476] = 33'b0100110000000000_1_0_xx_000_100_xxx_1_x_xx;
      patterns[5477] = 33'b0100110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5478] = 33'b0000010001011111_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5479] = 33'b0000110001011111_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5480] = 33'b0000110001011111_0_0_00_000_000_000_0_0_00;
      patterns[5481] = 33'b1000010000000101_0_1_00_000_101_100_0_x_00;
      patterns[5482] = 33'b1000110000000101_1_1_00_000_101_100_0_x_00;
      patterns[5483] = 33'b1000110000000101_0_0_00_000_000_000_0_0_00;
      patterns[5484] = 33'b1001010000000101_0_1_01_000_101_100_0_x_00;
      patterns[5485] = 33'b1001110000000101_1_1_01_000_101_100_0_x_00;
      patterns[5486] = 33'b1001110000000101_0_0_00_000_000_000_0_0_00;
      patterns[5487] = 33'b1010010000000101_0_1_10_000_101_100_0_x_00;
      patterns[5488] = 33'b1010110000000101_1_1_10_000_101_100_0_x_00;
      patterns[5489] = 33'b1010110000000101_0_0_00_000_000_000_0_0_00;
      patterns[5490] = 33'b1011010000000101_0_1_11_000_101_100_0_x_00;
      patterns[5491] = 33'b1011110000000101_1_1_11_000_101_100_0_x_00;
      patterns[5492] = 33'b1011110000000101_0_0_00_000_000_000_0_0_00;
      patterns[5493] = 33'b0101010000000000_0_1_xx_000_xxx_100_0_1_01;
      patterns[5494] = 33'b0101110000000000_1_1_xx_000_xxx_100_0_1_01;
      patterns[5495] = 33'b0101110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5496] = 33'b0100010000000000_0_0_xx_000_100_xxx_1_x_xx;
      patterns[5497] = 33'b0100110000000000_1_0_xx_000_100_xxx_1_x_xx;
      patterns[5498] = 33'b0100110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5499] = 33'b0000010011011111_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5500] = 33'b0000110011011111_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5501] = 33'b0000110011011111_0_0_00_000_000_000_0_0_00;
      patterns[5502] = 33'b1000010000000110_0_1_00_000_110_100_0_x_00;
      patterns[5503] = 33'b1000110000000110_1_1_00_000_110_100_0_x_00;
      patterns[5504] = 33'b1000110000000110_0_0_00_000_000_000_0_0_00;
      patterns[5505] = 33'b1001010000000110_0_1_01_000_110_100_0_x_00;
      patterns[5506] = 33'b1001110000000110_1_1_01_000_110_100_0_x_00;
      patterns[5507] = 33'b1001110000000110_0_0_00_000_000_000_0_0_00;
      patterns[5508] = 33'b1010010000000110_0_1_10_000_110_100_0_x_00;
      patterns[5509] = 33'b1010110000000110_1_1_10_000_110_100_0_x_00;
      patterns[5510] = 33'b1010110000000110_0_0_00_000_000_000_0_0_00;
      patterns[5511] = 33'b1011010000000110_0_1_11_000_110_100_0_x_00;
      patterns[5512] = 33'b1011110000000110_1_1_11_000_110_100_0_x_00;
      patterns[5513] = 33'b1011110000000110_0_0_00_000_000_000_0_0_00;
      patterns[5514] = 33'b0101010000000000_0_1_xx_000_xxx_100_0_1_01;
      patterns[5515] = 33'b0101110000000000_1_1_xx_000_xxx_100_0_1_01;
      patterns[5516] = 33'b0101110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5517] = 33'b0100010000000000_0_0_xx_000_100_xxx_1_x_xx;
      patterns[5518] = 33'b0100110000000000_1_0_xx_000_100_xxx_1_x_xx;
      patterns[5519] = 33'b0100110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5520] = 33'b0000010000110001_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5521] = 33'b0000110000110001_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5522] = 33'b0000110000110001_0_0_00_000_000_000_0_0_00;
      patterns[5523] = 33'b1000010000000111_0_1_00_000_111_100_0_x_00;
      patterns[5524] = 33'b1000110000000111_1_1_00_000_111_100_0_x_00;
      patterns[5525] = 33'b1000110000000111_0_0_00_000_000_000_0_0_00;
      patterns[5526] = 33'b1001010000000111_0_1_01_000_111_100_0_x_00;
      patterns[5527] = 33'b1001110000000111_1_1_01_000_111_100_0_x_00;
      patterns[5528] = 33'b1001110000000111_0_0_00_000_000_000_0_0_00;
      patterns[5529] = 33'b1010010000000111_0_1_10_000_111_100_0_x_00;
      patterns[5530] = 33'b1010110000000111_1_1_10_000_111_100_0_x_00;
      patterns[5531] = 33'b1010110000000111_0_0_00_000_000_000_0_0_00;
      patterns[5532] = 33'b1011010000000111_0_1_11_000_111_100_0_x_00;
      patterns[5533] = 33'b1011110000000111_1_1_11_000_111_100_0_x_00;
      patterns[5534] = 33'b1011110000000111_0_0_00_000_000_000_0_0_00;
      patterns[5535] = 33'b0101010000000000_0_1_xx_000_xxx_100_0_1_01;
      patterns[5536] = 33'b0101110000000000_1_1_xx_000_xxx_100_0_1_01;
      patterns[5537] = 33'b0101110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5538] = 33'b0100010000000000_0_0_xx_000_100_xxx_1_x_xx;
      patterns[5539] = 33'b0100110000000000_1_0_xx_000_100_xxx_1_x_xx;
      patterns[5540] = 33'b0100110000000000_0_0_00_000_000_000_0_0_00;
      patterns[5541] = 33'b0000010000010111_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5542] = 33'b0000110000010111_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5543] = 33'b0000110000010111_0_0_00_000_000_000_0_0_00;
      patterns[5544] = 33'b1000010000010000_0_1_00_001_000_100_0_x_00;
      patterns[5545] = 33'b1000110000010000_1_1_00_001_000_100_0_x_00;
      patterns[5546] = 33'b1000110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5547] = 33'b1001010000010000_0_1_01_001_000_100_0_x_00;
      patterns[5548] = 33'b1001110000010000_1_1_01_001_000_100_0_x_00;
      patterns[5549] = 33'b1001110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5550] = 33'b1010010000010000_0_1_10_001_000_100_0_x_00;
      patterns[5551] = 33'b1010110000010000_1_1_10_001_000_100_0_x_00;
      patterns[5552] = 33'b1010110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5553] = 33'b1011010000010000_0_1_11_001_000_100_0_x_00;
      patterns[5554] = 33'b1011110000010000_1_1_11_001_000_100_0_x_00;
      patterns[5555] = 33'b1011110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5556] = 33'b0101010000010000_0_1_xx_001_xxx_100_0_1_01;
      patterns[5557] = 33'b0101110000010000_1_1_xx_001_xxx_100_0_1_01;
      patterns[5558] = 33'b0101110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5559] = 33'b0100010000010000_0_0_xx_001_100_xxx_1_x_xx;
      patterns[5560] = 33'b0100110000010000_1_0_xx_001_100_xxx_1_x_xx;
      patterns[5561] = 33'b0100110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5562] = 33'b0000010011110110_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5563] = 33'b0000110011110110_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5564] = 33'b0000110011110110_0_0_00_000_000_000_0_0_00;
      patterns[5565] = 33'b1000010000010001_0_1_00_001_001_100_0_x_00;
      patterns[5566] = 33'b1000110000010001_1_1_00_001_001_100_0_x_00;
      patterns[5567] = 33'b1000110000010001_0_0_00_000_000_000_0_0_00;
      patterns[5568] = 33'b1001010000010001_0_1_01_001_001_100_0_x_00;
      patterns[5569] = 33'b1001110000010001_1_1_01_001_001_100_0_x_00;
      patterns[5570] = 33'b1001110000010001_0_0_00_000_000_000_0_0_00;
      patterns[5571] = 33'b1010010000010001_0_1_10_001_001_100_0_x_00;
      patterns[5572] = 33'b1010110000010001_1_1_10_001_001_100_0_x_00;
      patterns[5573] = 33'b1010110000010001_0_0_00_000_000_000_0_0_00;
      patterns[5574] = 33'b1011010000010001_0_1_11_001_001_100_0_x_00;
      patterns[5575] = 33'b1011110000010001_1_1_11_001_001_100_0_x_00;
      patterns[5576] = 33'b1011110000010001_0_0_00_000_000_000_0_0_00;
      patterns[5577] = 33'b0101010000010000_0_1_xx_001_xxx_100_0_1_01;
      patterns[5578] = 33'b0101110000010000_1_1_xx_001_xxx_100_0_1_01;
      patterns[5579] = 33'b0101110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5580] = 33'b0100010000010000_0_0_xx_001_100_xxx_1_x_xx;
      patterns[5581] = 33'b0100110000010000_1_0_xx_001_100_xxx_1_x_xx;
      patterns[5582] = 33'b0100110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5583] = 33'b0000010010111101_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5584] = 33'b0000110010111101_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5585] = 33'b0000110010111101_0_0_00_000_000_000_0_0_00;
      patterns[5586] = 33'b1000010000010010_0_1_00_001_010_100_0_x_00;
      patterns[5587] = 33'b1000110000010010_1_1_00_001_010_100_0_x_00;
      patterns[5588] = 33'b1000110000010010_0_0_00_000_000_000_0_0_00;
      patterns[5589] = 33'b1001010000010010_0_1_01_001_010_100_0_x_00;
      patterns[5590] = 33'b1001110000010010_1_1_01_001_010_100_0_x_00;
      patterns[5591] = 33'b1001110000010010_0_0_00_000_000_000_0_0_00;
      patterns[5592] = 33'b1010010000010010_0_1_10_001_010_100_0_x_00;
      patterns[5593] = 33'b1010110000010010_1_1_10_001_010_100_0_x_00;
      patterns[5594] = 33'b1010110000010010_0_0_00_000_000_000_0_0_00;
      patterns[5595] = 33'b1011010000010010_0_1_11_001_010_100_0_x_00;
      patterns[5596] = 33'b1011110000010010_1_1_11_001_010_100_0_x_00;
      patterns[5597] = 33'b1011110000010010_0_0_00_000_000_000_0_0_00;
      patterns[5598] = 33'b0101010000010000_0_1_xx_001_xxx_100_0_1_01;
      patterns[5599] = 33'b0101110000010000_1_1_xx_001_xxx_100_0_1_01;
      patterns[5600] = 33'b0101110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5601] = 33'b0100010000010000_0_0_xx_001_100_xxx_1_x_xx;
      patterns[5602] = 33'b0100110000010000_1_0_xx_001_100_xxx_1_x_xx;
      patterns[5603] = 33'b0100110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5604] = 33'b0000010010000111_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5605] = 33'b0000110010000111_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5606] = 33'b0000110010000111_0_0_00_000_000_000_0_0_00;
      patterns[5607] = 33'b1000010000010011_0_1_00_001_011_100_0_x_00;
      patterns[5608] = 33'b1000110000010011_1_1_00_001_011_100_0_x_00;
      patterns[5609] = 33'b1000110000010011_0_0_00_000_000_000_0_0_00;
      patterns[5610] = 33'b1001010000010011_0_1_01_001_011_100_0_x_00;
      patterns[5611] = 33'b1001110000010011_1_1_01_001_011_100_0_x_00;
      patterns[5612] = 33'b1001110000010011_0_0_00_000_000_000_0_0_00;
      patterns[5613] = 33'b1010010000010011_0_1_10_001_011_100_0_x_00;
      patterns[5614] = 33'b1010110000010011_1_1_10_001_011_100_0_x_00;
      patterns[5615] = 33'b1010110000010011_0_0_00_000_000_000_0_0_00;
      patterns[5616] = 33'b1011010000010011_0_1_11_001_011_100_0_x_00;
      patterns[5617] = 33'b1011110000010011_1_1_11_001_011_100_0_x_00;
      patterns[5618] = 33'b1011110000010011_0_0_00_000_000_000_0_0_00;
      patterns[5619] = 33'b0101010000010000_0_1_xx_001_xxx_100_0_1_01;
      patterns[5620] = 33'b0101110000010000_1_1_xx_001_xxx_100_0_1_01;
      patterns[5621] = 33'b0101110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5622] = 33'b0100010000010000_0_0_xx_001_100_xxx_1_x_xx;
      patterns[5623] = 33'b0100110000010000_1_0_xx_001_100_xxx_1_x_xx;
      patterns[5624] = 33'b0100110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5625] = 33'b0000010001100110_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5626] = 33'b0000110001100110_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5627] = 33'b0000110001100110_0_0_00_000_000_000_0_0_00;
      patterns[5628] = 33'b1000010000010100_0_1_00_001_100_100_0_x_00;
      patterns[5629] = 33'b1000110000010100_1_1_00_001_100_100_0_x_00;
      patterns[5630] = 33'b1000110000010100_0_0_00_000_000_000_0_0_00;
      patterns[5631] = 33'b1001010000010100_0_1_01_001_100_100_0_x_00;
      patterns[5632] = 33'b1001110000010100_1_1_01_001_100_100_0_x_00;
      patterns[5633] = 33'b1001110000010100_0_0_00_000_000_000_0_0_00;
      patterns[5634] = 33'b1010010000010100_0_1_10_001_100_100_0_x_00;
      patterns[5635] = 33'b1010110000010100_1_1_10_001_100_100_0_x_00;
      patterns[5636] = 33'b1010110000010100_0_0_00_000_000_000_0_0_00;
      patterns[5637] = 33'b1011010000010100_0_1_11_001_100_100_0_x_00;
      patterns[5638] = 33'b1011110000010100_1_1_11_001_100_100_0_x_00;
      patterns[5639] = 33'b1011110000010100_0_0_00_000_000_000_0_0_00;
      patterns[5640] = 33'b0101010000010000_0_1_xx_001_xxx_100_0_1_01;
      patterns[5641] = 33'b0101110000010000_1_1_xx_001_xxx_100_0_1_01;
      patterns[5642] = 33'b0101110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5643] = 33'b0100010000010000_0_0_xx_001_100_xxx_1_x_xx;
      patterns[5644] = 33'b0100110000010000_1_0_xx_001_100_xxx_1_x_xx;
      patterns[5645] = 33'b0100110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5646] = 33'b0000010000101000_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5647] = 33'b0000110000101000_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5648] = 33'b0000110000101000_0_0_00_000_000_000_0_0_00;
      patterns[5649] = 33'b1000010000010101_0_1_00_001_101_100_0_x_00;
      patterns[5650] = 33'b1000110000010101_1_1_00_001_101_100_0_x_00;
      patterns[5651] = 33'b1000110000010101_0_0_00_000_000_000_0_0_00;
      patterns[5652] = 33'b1001010000010101_0_1_01_001_101_100_0_x_00;
      patterns[5653] = 33'b1001110000010101_1_1_01_001_101_100_0_x_00;
      patterns[5654] = 33'b1001110000010101_0_0_00_000_000_000_0_0_00;
      patterns[5655] = 33'b1010010000010101_0_1_10_001_101_100_0_x_00;
      patterns[5656] = 33'b1010110000010101_1_1_10_001_101_100_0_x_00;
      patterns[5657] = 33'b1010110000010101_0_0_00_000_000_000_0_0_00;
      patterns[5658] = 33'b1011010000010101_0_1_11_001_101_100_0_x_00;
      patterns[5659] = 33'b1011110000010101_1_1_11_001_101_100_0_x_00;
      patterns[5660] = 33'b1011110000010101_0_0_00_000_000_000_0_0_00;
      patterns[5661] = 33'b0101010000010000_0_1_xx_001_xxx_100_0_1_01;
      patterns[5662] = 33'b0101110000010000_1_1_xx_001_xxx_100_0_1_01;
      patterns[5663] = 33'b0101110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5664] = 33'b0100010000010000_0_0_xx_001_100_xxx_1_x_xx;
      patterns[5665] = 33'b0100110000010000_1_0_xx_001_100_xxx_1_x_xx;
      patterns[5666] = 33'b0100110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5667] = 33'b0000010001100010_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5668] = 33'b0000110001100010_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5669] = 33'b0000110001100010_0_0_00_000_000_000_0_0_00;
      patterns[5670] = 33'b1000010000010110_0_1_00_001_110_100_0_x_00;
      patterns[5671] = 33'b1000110000010110_1_1_00_001_110_100_0_x_00;
      patterns[5672] = 33'b1000110000010110_0_0_00_000_000_000_0_0_00;
      patterns[5673] = 33'b1001010000010110_0_1_01_001_110_100_0_x_00;
      patterns[5674] = 33'b1001110000010110_1_1_01_001_110_100_0_x_00;
      patterns[5675] = 33'b1001110000010110_0_0_00_000_000_000_0_0_00;
      patterns[5676] = 33'b1010010000010110_0_1_10_001_110_100_0_x_00;
      patterns[5677] = 33'b1010110000010110_1_1_10_001_110_100_0_x_00;
      patterns[5678] = 33'b1010110000010110_0_0_00_000_000_000_0_0_00;
      patterns[5679] = 33'b1011010000010110_0_1_11_001_110_100_0_x_00;
      patterns[5680] = 33'b1011110000010110_1_1_11_001_110_100_0_x_00;
      patterns[5681] = 33'b1011110000010110_0_0_00_000_000_000_0_0_00;
      patterns[5682] = 33'b0101010000010000_0_1_xx_001_xxx_100_0_1_01;
      patterns[5683] = 33'b0101110000010000_1_1_xx_001_xxx_100_0_1_01;
      patterns[5684] = 33'b0101110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5685] = 33'b0100010000010000_0_0_xx_001_100_xxx_1_x_xx;
      patterns[5686] = 33'b0100110000010000_1_0_xx_001_100_xxx_1_x_xx;
      patterns[5687] = 33'b0100110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5688] = 33'b0000010011100001_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5689] = 33'b0000110011100001_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5690] = 33'b0000110011100001_0_0_00_000_000_000_0_0_00;
      patterns[5691] = 33'b1000010000010111_0_1_00_001_111_100_0_x_00;
      patterns[5692] = 33'b1000110000010111_1_1_00_001_111_100_0_x_00;
      patterns[5693] = 33'b1000110000010111_0_0_00_000_000_000_0_0_00;
      patterns[5694] = 33'b1001010000010111_0_1_01_001_111_100_0_x_00;
      patterns[5695] = 33'b1001110000010111_1_1_01_001_111_100_0_x_00;
      patterns[5696] = 33'b1001110000010111_0_0_00_000_000_000_0_0_00;
      patterns[5697] = 33'b1010010000010111_0_1_10_001_111_100_0_x_00;
      patterns[5698] = 33'b1010110000010111_1_1_10_001_111_100_0_x_00;
      patterns[5699] = 33'b1010110000010111_0_0_00_000_000_000_0_0_00;
      patterns[5700] = 33'b1011010000010111_0_1_11_001_111_100_0_x_00;
      patterns[5701] = 33'b1011110000010111_1_1_11_001_111_100_0_x_00;
      patterns[5702] = 33'b1011110000010111_0_0_00_000_000_000_0_0_00;
      patterns[5703] = 33'b0101010000010000_0_1_xx_001_xxx_100_0_1_01;
      patterns[5704] = 33'b0101110000010000_1_1_xx_001_xxx_100_0_1_01;
      patterns[5705] = 33'b0101110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5706] = 33'b0100010000010000_0_0_xx_001_100_xxx_1_x_xx;
      patterns[5707] = 33'b0100110000010000_1_0_xx_001_100_xxx_1_x_xx;
      patterns[5708] = 33'b0100110000010000_0_0_00_000_000_000_0_0_00;
      patterns[5709] = 33'b0000010011011110_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5710] = 33'b0000110011011110_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5711] = 33'b0000110011011110_0_0_00_000_000_000_0_0_00;
      patterns[5712] = 33'b1000010000100000_0_1_00_010_000_100_0_x_00;
      patterns[5713] = 33'b1000110000100000_1_1_00_010_000_100_0_x_00;
      patterns[5714] = 33'b1000110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5715] = 33'b1001010000100000_0_1_01_010_000_100_0_x_00;
      patterns[5716] = 33'b1001110000100000_1_1_01_010_000_100_0_x_00;
      patterns[5717] = 33'b1001110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5718] = 33'b1010010000100000_0_1_10_010_000_100_0_x_00;
      patterns[5719] = 33'b1010110000100000_1_1_10_010_000_100_0_x_00;
      patterns[5720] = 33'b1010110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5721] = 33'b1011010000100000_0_1_11_010_000_100_0_x_00;
      patterns[5722] = 33'b1011110000100000_1_1_11_010_000_100_0_x_00;
      patterns[5723] = 33'b1011110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5724] = 33'b0101010000100000_0_1_xx_010_xxx_100_0_1_01;
      patterns[5725] = 33'b0101110000100000_1_1_xx_010_xxx_100_0_1_01;
      patterns[5726] = 33'b0101110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5727] = 33'b0100010000100000_0_0_xx_010_100_xxx_1_x_xx;
      patterns[5728] = 33'b0100110000100000_1_0_xx_010_100_xxx_1_x_xx;
      patterns[5729] = 33'b0100110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5730] = 33'b0000010001000110_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5731] = 33'b0000110001000110_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5732] = 33'b0000110001000110_0_0_00_000_000_000_0_0_00;
      patterns[5733] = 33'b1000010000100001_0_1_00_010_001_100_0_x_00;
      patterns[5734] = 33'b1000110000100001_1_1_00_010_001_100_0_x_00;
      patterns[5735] = 33'b1000110000100001_0_0_00_000_000_000_0_0_00;
      patterns[5736] = 33'b1001010000100001_0_1_01_010_001_100_0_x_00;
      patterns[5737] = 33'b1001110000100001_1_1_01_010_001_100_0_x_00;
      patterns[5738] = 33'b1001110000100001_0_0_00_000_000_000_0_0_00;
      patterns[5739] = 33'b1010010000100001_0_1_10_010_001_100_0_x_00;
      patterns[5740] = 33'b1010110000100001_1_1_10_010_001_100_0_x_00;
      patterns[5741] = 33'b1010110000100001_0_0_00_000_000_000_0_0_00;
      patterns[5742] = 33'b1011010000100001_0_1_11_010_001_100_0_x_00;
      patterns[5743] = 33'b1011110000100001_1_1_11_010_001_100_0_x_00;
      patterns[5744] = 33'b1011110000100001_0_0_00_000_000_000_0_0_00;
      patterns[5745] = 33'b0101010000100000_0_1_xx_010_xxx_100_0_1_01;
      patterns[5746] = 33'b0101110000100000_1_1_xx_010_xxx_100_0_1_01;
      patterns[5747] = 33'b0101110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5748] = 33'b0100010000100000_0_0_xx_010_100_xxx_1_x_xx;
      patterns[5749] = 33'b0100110000100000_1_0_xx_010_100_xxx_1_x_xx;
      patterns[5750] = 33'b0100110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5751] = 33'b0000010000110011_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5752] = 33'b0000110000110011_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5753] = 33'b0000110000110011_0_0_00_000_000_000_0_0_00;
      patterns[5754] = 33'b1000010000100010_0_1_00_010_010_100_0_x_00;
      patterns[5755] = 33'b1000110000100010_1_1_00_010_010_100_0_x_00;
      patterns[5756] = 33'b1000110000100010_0_0_00_000_000_000_0_0_00;
      patterns[5757] = 33'b1001010000100010_0_1_01_010_010_100_0_x_00;
      patterns[5758] = 33'b1001110000100010_1_1_01_010_010_100_0_x_00;
      patterns[5759] = 33'b1001110000100010_0_0_00_000_000_000_0_0_00;
      patterns[5760] = 33'b1010010000100010_0_1_10_010_010_100_0_x_00;
      patterns[5761] = 33'b1010110000100010_1_1_10_010_010_100_0_x_00;
      patterns[5762] = 33'b1010110000100010_0_0_00_000_000_000_0_0_00;
      patterns[5763] = 33'b1011010000100010_0_1_11_010_010_100_0_x_00;
      patterns[5764] = 33'b1011110000100010_1_1_11_010_010_100_0_x_00;
      patterns[5765] = 33'b1011110000100010_0_0_00_000_000_000_0_0_00;
      patterns[5766] = 33'b0101010000100000_0_1_xx_010_xxx_100_0_1_01;
      patterns[5767] = 33'b0101110000100000_1_1_xx_010_xxx_100_0_1_01;
      patterns[5768] = 33'b0101110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5769] = 33'b0100010000100000_0_0_xx_010_100_xxx_1_x_xx;
      patterns[5770] = 33'b0100110000100000_1_0_xx_010_100_xxx_1_x_xx;
      patterns[5771] = 33'b0100110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5772] = 33'b0000010000000101_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5773] = 33'b0000110000000101_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5774] = 33'b0000110000000101_0_0_00_000_000_000_0_0_00;
      patterns[5775] = 33'b1000010000100011_0_1_00_010_011_100_0_x_00;
      patterns[5776] = 33'b1000110000100011_1_1_00_010_011_100_0_x_00;
      patterns[5777] = 33'b1000110000100011_0_0_00_000_000_000_0_0_00;
      patterns[5778] = 33'b1001010000100011_0_1_01_010_011_100_0_x_00;
      patterns[5779] = 33'b1001110000100011_1_1_01_010_011_100_0_x_00;
      patterns[5780] = 33'b1001110000100011_0_0_00_000_000_000_0_0_00;
      patterns[5781] = 33'b1010010000100011_0_1_10_010_011_100_0_x_00;
      patterns[5782] = 33'b1010110000100011_1_1_10_010_011_100_0_x_00;
      patterns[5783] = 33'b1010110000100011_0_0_00_000_000_000_0_0_00;
      patterns[5784] = 33'b1011010000100011_0_1_11_010_011_100_0_x_00;
      patterns[5785] = 33'b1011110000100011_1_1_11_010_011_100_0_x_00;
      patterns[5786] = 33'b1011110000100011_0_0_00_000_000_000_0_0_00;
      patterns[5787] = 33'b0101010000100000_0_1_xx_010_xxx_100_0_1_01;
      patterns[5788] = 33'b0101110000100000_1_1_xx_010_xxx_100_0_1_01;
      patterns[5789] = 33'b0101110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5790] = 33'b0100010000100000_0_0_xx_010_100_xxx_1_x_xx;
      patterns[5791] = 33'b0100110000100000_1_0_xx_010_100_xxx_1_x_xx;
      patterns[5792] = 33'b0100110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5793] = 33'b0000010000111001_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5794] = 33'b0000110000111001_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5795] = 33'b0000110000111001_0_0_00_000_000_000_0_0_00;
      patterns[5796] = 33'b1000010000100100_0_1_00_010_100_100_0_x_00;
      patterns[5797] = 33'b1000110000100100_1_1_00_010_100_100_0_x_00;
      patterns[5798] = 33'b1000110000100100_0_0_00_000_000_000_0_0_00;
      patterns[5799] = 33'b1001010000100100_0_1_01_010_100_100_0_x_00;
      patterns[5800] = 33'b1001110000100100_1_1_01_010_100_100_0_x_00;
      patterns[5801] = 33'b1001110000100100_0_0_00_000_000_000_0_0_00;
      patterns[5802] = 33'b1010010000100100_0_1_10_010_100_100_0_x_00;
      patterns[5803] = 33'b1010110000100100_1_1_10_010_100_100_0_x_00;
      patterns[5804] = 33'b1010110000100100_0_0_00_000_000_000_0_0_00;
      patterns[5805] = 33'b1011010000100100_0_1_11_010_100_100_0_x_00;
      patterns[5806] = 33'b1011110000100100_1_1_11_010_100_100_0_x_00;
      patterns[5807] = 33'b1011110000100100_0_0_00_000_000_000_0_0_00;
      patterns[5808] = 33'b0101010000100000_0_1_xx_010_xxx_100_0_1_01;
      patterns[5809] = 33'b0101110000100000_1_1_xx_010_xxx_100_0_1_01;
      patterns[5810] = 33'b0101110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5811] = 33'b0100010000100000_0_0_xx_010_100_xxx_1_x_xx;
      patterns[5812] = 33'b0100110000100000_1_0_xx_010_100_xxx_1_x_xx;
      patterns[5813] = 33'b0100110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5814] = 33'b0000010001101001_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5815] = 33'b0000110001101001_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5816] = 33'b0000110001101001_0_0_00_000_000_000_0_0_00;
      patterns[5817] = 33'b1000010000100101_0_1_00_010_101_100_0_x_00;
      patterns[5818] = 33'b1000110000100101_1_1_00_010_101_100_0_x_00;
      patterns[5819] = 33'b1000110000100101_0_0_00_000_000_000_0_0_00;
      patterns[5820] = 33'b1001010000100101_0_1_01_010_101_100_0_x_00;
      patterns[5821] = 33'b1001110000100101_1_1_01_010_101_100_0_x_00;
      patterns[5822] = 33'b1001110000100101_0_0_00_000_000_000_0_0_00;
      patterns[5823] = 33'b1010010000100101_0_1_10_010_101_100_0_x_00;
      patterns[5824] = 33'b1010110000100101_1_1_10_010_101_100_0_x_00;
      patterns[5825] = 33'b1010110000100101_0_0_00_000_000_000_0_0_00;
      patterns[5826] = 33'b1011010000100101_0_1_11_010_101_100_0_x_00;
      patterns[5827] = 33'b1011110000100101_1_1_11_010_101_100_0_x_00;
      patterns[5828] = 33'b1011110000100101_0_0_00_000_000_000_0_0_00;
      patterns[5829] = 33'b0101010000100000_0_1_xx_010_xxx_100_0_1_01;
      patterns[5830] = 33'b0101110000100000_1_1_xx_010_xxx_100_0_1_01;
      patterns[5831] = 33'b0101110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5832] = 33'b0100010000100000_0_0_xx_010_100_xxx_1_x_xx;
      patterns[5833] = 33'b0100110000100000_1_0_xx_010_100_xxx_1_x_xx;
      patterns[5834] = 33'b0100110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5835] = 33'b0000010011011110_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5836] = 33'b0000110011011110_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5837] = 33'b0000110011011110_0_0_00_000_000_000_0_0_00;
      patterns[5838] = 33'b1000010000100110_0_1_00_010_110_100_0_x_00;
      patterns[5839] = 33'b1000110000100110_1_1_00_010_110_100_0_x_00;
      patterns[5840] = 33'b1000110000100110_0_0_00_000_000_000_0_0_00;
      patterns[5841] = 33'b1001010000100110_0_1_01_010_110_100_0_x_00;
      patterns[5842] = 33'b1001110000100110_1_1_01_010_110_100_0_x_00;
      patterns[5843] = 33'b1001110000100110_0_0_00_000_000_000_0_0_00;
      patterns[5844] = 33'b1010010000100110_0_1_10_010_110_100_0_x_00;
      patterns[5845] = 33'b1010110000100110_1_1_10_010_110_100_0_x_00;
      patterns[5846] = 33'b1010110000100110_0_0_00_000_000_000_0_0_00;
      patterns[5847] = 33'b1011010000100110_0_1_11_010_110_100_0_x_00;
      patterns[5848] = 33'b1011110000100110_1_1_11_010_110_100_0_x_00;
      patterns[5849] = 33'b1011110000100110_0_0_00_000_000_000_0_0_00;
      patterns[5850] = 33'b0101010000100000_0_1_xx_010_xxx_100_0_1_01;
      patterns[5851] = 33'b0101110000100000_1_1_xx_010_xxx_100_0_1_01;
      patterns[5852] = 33'b0101110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5853] = 33'b0100010000100000_0_0_xx_010_100_xxx_1_x_xx;
      patterns[5854] = 33'b0100110000100000_1_0_xx_010_100_xxx_1_x_xx;
      patterns[5855] = 33'b0100110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5856] = 33'b0000010011101001_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5857] = 33'b0000110011101001_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5858] = 33'b0000110011101001_0_0_00_000_000_000_0_0_00;
      patterns[5859] = 33'b1000010000100111_0_1_00_010_111_100_0_x_00;
      patterns[5860] = 33'b1000110000100111_1_1_00_010_111_100_0_x_00;
      patterns[5861] = 33'b1000110000100111_0_0_00_000_000_000_0_0_00;
      patterns[5862] = 33'b1001010000100111_0_1_01_010_111_100_0_x_00;
      patterns[5863] = 33'b1001110000100111_1_1_01_010_111_100_0_x_00;
      patterns[5864] = 33'b1001110000100111_0_0_00_000_000_000_0_0_00;
      patterns[5865] = 33'b1010010000100111_0_1_10_010_111_100_0_x_00;
      patterns[5866] = 33'b1010110000100111_1_1_10_010_111_100_0_x_00;
      patterns[5867] = 33'b1010110000100111_0_0_00_000_000_000_0_0_00;
      patterns[5868] = 33'b1011010000100111_0_1_11_010_111_100_0_x_00;
      patterns[5869] = 33'b1011110000100111_1_1_11_010_111_100_0_x_00;
      patterns[5870] = 33'b1011110000100111_0_0_00_000_000_000_0_0_00;
      patterns[5871] = 33'b0101010000100000_0_1_xx_010_xxx_100_0_1_01;
      patterns[5872] = 33'b0101110000100000_1_1_xx_010_xxx_100_0_1_01;
      patterns[5873] = 33'b0101110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5874] = 33'b0100010000100000_0_0_xx_010_100_xxx_1_x_xx;
      patterns[5875] = 33'b0100110000100000_1_0_xx_010_100_xxx_1_x_xx;
      patterns[5876] = 33'b0100110000100000_0_0_00_000_000_000_0_0_00;
      patterns[5877] = 33'b0000010011001001_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5878] = 33'b0000110011001001_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5879] = 33'b0000110011001001_0_0_00_000_000_000_0_0_00;
      patterns[5880] = 33'b1000010000110000_0_1_00_011_000_100_0_x_00;
      patterns[5881] = 33'b1000110000110000_1_1_00_011_000_100_0_x_00;
      patterns[5882] = 33'b1000110000110000_0_0_00_000_000_000_0_0_00;
      patterns[5883] = 33'b1001010000110000_0_1_01_011_000_100_0_x_00;
      patterns[5884] = 33'b1001110000110000_1_1_01_011_000_100_0_x_00;
      patterns[5885] = 33'b1001110000110000_0_0_00_000_000_000_0_0_00;
      patterns[5886] = 33'b1010010000110000_0_1_10_011_000_100_0_x_00;
      patterns[5887] = 33'b1010110000110000_1_1_10_011_000_100_0_x_00;
      patterns[5888] = 33'b1010110000110000_0_0_00_000_000_000_0_0_00;
      patterns[5889] = 33'b1011010000110000_0_1_11_011_000_100_0_x_00;
      patterns[5890] = 33'b1011110000110000_1_1_11_011_000_100_0_x_00;
      patterns[5891] = 33'b1011110000110000_0_0_00_000_000_000_0_0_00;
      patterns[5892] = 33'b0101010000110000_0_1_xx_011_xxx_100_0_1_01;
      patterns[5893] = 33'b0101110000110000_1_1_xx_011_xxx_100_0_1_01;
      patterns[5894] = 33'b0101110000110000_0_0_00_000_000_000_0_0_00;
      patterns[5895] = 33'b0100010000110000_0_0_xx_011_100_xxx_1_x_xx;
      patterns[5896] = 33'b0100110000110000_1_0_xx_011_100_xxx_1_x_xx;
      patterns[5897] = 33'b0100110000110000_0_0_00_000_000_000_0_0_00;
      patterns[5898] = 33'b0000010001110111_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5899] = 33'b0000110001110111_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5900] = 33'b0000110001110111_0_0_00_000_000_000_0_0_00;
      patterns[5901] = 33'b1000010000110001_0_1_00_011_001_100_0_x_00;
      patterns[5902] = 33'b1000110000110001_1_1_00_011_001_100_0_x_00;
      patterns[5903] = 33'b1000110000110001_0_0_00_000_000_000_0_0_00;
      patterns[5904] = 33'b1001010000110001_0_1_01_011_001_100_0_x_00;
      patterns[5905] = 33'b1001110000110001_1_1_01_011_001_100_0_x_00;
      patterns[5906] = 33'b1001110000110001_0_0_00_000_000_000_0_0_00;
      patterns[5907] = 33'b1010010000110001_0_1_10_011_001_100_0_x_00;
      patterns[5908] = 33'b1010110000110001_1_1_10_011_001_100_0_x_00;
      patterns[5909] = 33'b1010110000110001_0_0_00_000_000_000_0_0_00;
      patterns[5910] = 33'b1011010000110001_0_1_11_011_001_100_0_x_00;
      patterns[5911] = 33'b1011110000110001_1_1_11_011_001_100_0_x_00;
      patterns[5912] = 33'b1011110000110001_0_0_00_000_000_000_0_0_00;
      patterns[5913] = 33'b0101010000110000_0_1_xx_011_xxx_100_0_1_01;
      patterns[5914] = 33'b0101110000110000_1_1_xx_011_xxx_100_0_1_01;
      patterns[5915] = 33'b0101110000110000_0_0_00_000_000_000_0_0_00;
      patterns[5916] = 33'b0100010000110000_0_0_xx_011_100_xxx_1_x_xx;
      patterns[5917] = 33'b0100110000110000_1_0_xx_011_100_xxx_1_x_xx;
      patterns[5918] = 33'b0100110000110000_0_0_00_000_000_000_0_0_00;
      patterns[5919] = 33'b0000010011101011_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5920] = 33'b0000110011101011_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5921] = 33'b0000110011101011_0_0_00_000_000_000_0_0_00;
      patterns[5922] = 33'b1000010000110010_0_1_00_011_010_100_0_x_00;
      patterns[5923] = 33'b1000110000110010_1_1_00_011_010_100_0_x_00;
      patterns[5924] = 33'b1000110000110010_0_0_00_000_000_000_0_0_00;
      patterns[5925] = 33'b1001010000110010_0_1_01_011_010_100_0_x_00;
      patterns[5926] = 33'b1001110000110010_1_1_01_011_010_100_0_x_00;
      patterns[5927] = 33'b1001110000110010_0_0_00_000_000_000_0_0_00;
      patterns[5928] = 33'b1010010000110010_0_1_10_011_010_100_0_x_00;
      patterns[5929] = 33'b1010110000110010_1_1_10_011_010_100_0_x_00;
      patterns[5930] = 33'b1010110000110010_0_0_00_000_000_000_0_0_00;
      patterns[5931] = 33'b1011010000110010_0_1_11_011_010_100_0_x_00;
      patterns[5932] = 33'b1011110000110010_1_1_11_011_010_100_0_x_00;
      patterns[5933] = 33'b1011110000110010_0_0_00_000_000_000_0_0_00;
      patterns[5934] = 33'b0101010000110000_0_1_xx_011_xxx_100_0_1_01;
      patterns[5935] = 33'b0101110000110000_1_1_xx_011_xxx_100_0_1_01;
      patterns[5936] = 33'b0101110000110000_0_0_00_000_000_000_0_0_00;
      patterns[5937] = 33'b0100010000110000_0_0_xx_011_100_xxx_1_x_xx;
      patterns[5938] = 33'b0100110000110000_1_0_xx_011_100_xxx_1_x_xx;
      patterns[5939] = 33'b0100110000110000_0_0_00_000_000_000_0_0_00;
      patterns[5940] = 33'b0000010010101001_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5941] = 33'b0000110010101001_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5942] = 33'b0000110010101001_0_0_00_000_000_000_0_0_00;
      patterns[5943] = 33'b1000010000110011_0_1_00_011_011_100_0_x_00;
      patterns[5944] = 33'b1000110000110011_1_1_00_011_011_100_0_x_00;
      patterns[5945] = 33'b1000110000110011_0_0_00_000_000_000_0_0_00;
      patterns[5946] = 33'b1001010000110011_0_1_01_011_011_100_0_x_00;
      patterns[5947] = 33'b1001110000110011_1_1_01_011_011_100_0_x_00;
      patterns[5948] = 33'b1001110000110011_0_0_00_000_000_000_0_0_00;
      patterns[5949] = 33'b1010010000110011_0_1_10_011_011_100_0_x_00;
      patterns[5950] = 33'b1010110000110011_1_1_10_011_011_100_0_x_00;
      patterns[5951] = 33'b1010110000110011_0_0_00_000_000_000_0_0_00;
      patterns[5952] = 33'b1011010000110011_0_1_11_011_011_100_0_x_00;
      patterns[5953] = 33'b1011110000110011_1_1_11_011_011_100_0_x_00;
      patterns[5954] = 33'b1011110000110011_0_0_00_000_000_000_0_0_00;
      patterns[5955] = 33'b0101010000110000_0_1_xx_011_xxx_100_0_1_01;
      patterns[5956] = 33'b0101110000110000_1_1_xx_011_xxx_100_0_1_01;
      patterns[5957] = 33'b0101110000110000_0_0_00_000_000_000_0_0_00;
      patterns[5958] = 33'b0100010000110000_0_0_xx_011_100_xxx_1_x_xx;
      patterns[5959] = 33'b0100110000110000_1_0_xx_011_100_xxx_1_x_xx;
      patterns[5960] = 33'b0100110000110000_0_0_00_000_000_000_0_0_00;
      patterns[5961] = 33'b0000010010110111_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5962] = 33'b0000110010110111_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5963] = 33'b0000110010110111_0_0_00_000_000_000_0_0_00;
      patterns[5964] = 33'b1000010000110100_0_1_00_011_100_100_0_x_00;
      patterns[5965] = 33'b1000110000110100_1_1_00_011_100_100_0_x_00;
      patterns[5966] = 33'b1000110000110100_0_0_00_000_000_000_0_0_00;
      patterns[5967] = 33'b1001010000110100_0_1_01_011_100_100_0_x_00;
      patterns[5968] = 33'b1001110000110100_1_1_01_011_100_100_0_x_00;
      patterns[5969] = 33'b1001110000110100_0_0_00_000_000_000_0_0_00;
      patterns[5970] = 33'b1010010000110100_0_1_10_011_100_100_0_x_00;
      patterns[5971] = 33'b1010110000110100_1_1_10_011_100_100_0_x_00;
      patterns[5972] = 33'b1010110000110100_0_0_00_000_000_000_0_0_00;
      patterns[5973] = 33'b1011010000110100_0_1_11_011_100_100_0_x_00;
      patterns[5974] = 33'b1011110000110100_1_1_11_011_100_100_0_x_00;
      patterns[5975] = 33'b1011110000110100_0_0_00_000_000_000_0_0_00;
      patterns[5976] = 33'b0101010000110000_0_1_xx_011_xxx_100_0_1_01;
      patterns[5977] = 33'b0101110000110000_1_1_xx_011_xxx_100_0_1_01;
      patterns[5978] = 33'b0101110000110000_0_0_00_000_000_000_0_0_00;
      patterns[5979] = 33'b0100010000110000_0_0_xx_011_100_xxx_1_x_xx;
      patterns[5980] = 33'b0100110000110000_1_0_xx_011_100_xxx_1_x_xx;
      patterns[5981] = 33'b0100110000110000_0_0_00_000_000_000_0_0_00;
      patterns[5982] = 33'b0000010011111000_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[5983] = 33'b0000110011111000_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[5984] = 33'b0000110011111000_0_0_00_000_000_000_0_0_00;
      patterns[5985] = 33'b1000010000110101_0_1_00_011_101_100_0_x_00;
      patterns[5986] = 33'b1000110000110101_1_1_00_011_101_100_0_x_00;
      patterns[5987] = 33'b1000110000110101_0_0_00_000_000_000_0_0_00;
      patterns[5988] = 33'b1001010000110101_0_1_01_011_101_100_0_x_00;
      patterns[5989] = 33'b1001110000110101_1_1_01_011_101_100_0_x_00;
      patterns[5990] = 33'b1001110000110101_0_0_00_000_000_000_0_0_00;
      patterns[5991] = 33'b1010010000110101_0_1_10_011_101_100_0_x_00;
      patterns[5992] = 33'b1010110000110101_1_1_10_011_101_100_0_x_00;
      patterns[5993] = 33'b1010110000110101_0_0_00_000_000_000_0_0_00;
      patterns[5994] = 33'b1011010000110101_0_1_11_011_101_100_0_x_00;
      patterns[5995] = 33'b1011110000110101_1_1_11_011_101_100_0_x_00;
      patterns[5996] = 33'b1011110000110101_0_0_00_000_000_000_0_0_00;
      patterns[5997] = 33'b0101010000110000_0_1_xx_011_xxx_100_0_1_01;
      patterns[5998] = 33'b0101110000110000_1_1_xx_011_xxx_100_0_1_01;
      patterns[5999] = 33'b0101110000110000_0_0_00_000_000_000_0_0_00;
      patterns[6000] = 33'b0100010000110000_0_0_xx_011_100_xxx_1_x_xx;
      patterns[6001] = 33'b0100110000110000_1_0_xx_011_100_xxx_1_x_xx;
      patterns[6002] = 33'b0100110000110000_0_0_00_000_000_000_0_0_00;
      patterns[6003] = 33'b0000010010111011_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6004] = 33'b0000110010111011_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6005] = 33'b0000110010111011_0_0_00_000_000_000_0_0_00;
      patterns[6006] = 33'b1000010000110110_0_1_00_011_110_100_0_x_00;
      patterns[6007] = 33'b1000110000110110_1_1_00_011_110_100_0_x_00;
      patterns[6008] = 33'b1000110000110110_0_0_00_000_000_000_0_0_00;
      patterns[6009] = 33'b1001010000110110_0_1_01_011_110_100_0_x_00;
      patterns[6010] = 33'b1001110000110110_1_1_01_011_110_100_0_x_00;
      patterns[6011] = 33'b1001110000110110_0_0_00_000_000_000_0_0_00;
      patterns[6012] = 33'b1010010000110110_0_1_10_011_110_100_0_x_00;
      patterns[6013] = 33'b1010110000110110_1_1_10_011_110_100_0_x_00;
      patterns[6014] = 33'b1010110000110110_0_0_00_000_000_000_0_0_00;
      patterns[6015] = 33'b1011010000110110_0_1_11_011_110_100_0_x_00;
      patterns[6016] = 33'b1011110000110110_1_1_11_011_110_100_0_x_00;
      patterns[6017] = 33'b1011110000110110_0_0_00_000_000_000_0_0_00;
      patterns[6018] = 33'b0101010000110000_0_1_xx_011_xxx_100_0_1_01;
      patterns[6019] = 33'b0101110000110000_1_1_xx_011_xxx_100_0_1_01;
      patterns[6020] = 33'b0101110000110000_0_0_00_000_000_000_0_0_00;
      patterns[6021] = 33'b0100010000110000_0_0_xx_011_100_xxx_1_x_xx;
      patterns[6022] = 33'b0100110000110000_1_0_xx_011_100_xxx_1_x_xx;
      patterns[6023] = 33'b0100110000110000_0_0_00_000_000_000_0_0_00;
      patterns[6024] = 33'b0000010000100101_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6025] = 33'b0000110000100101_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6026] = 33'b0000110000100101_0_0_00_000_000_000_0_0_00;
      patterns[6027] = 33'b1000010000110111_0_1_00_011_111_100_0_x_00;
      patterns[6028] = 33'b1000110000110111_1_1_00_011_111_100_0_x_00;
      patterns[6029] = 33'b1000110000110111_0_0_00_000_000_000_0_0_00;
      patterns[6030] = 33'b1001010000110111_0_1_01_011_111_100_0_x_00;
      patterns[6031] = 33'b1001110000110111_1_1_01_011_111_100_0_x_00;
      patterns[6032] = 33'b1001110000110111_0_0_00_000_000_000_0_0_00;
      patterns[6033] = 33'b1010010000110111_0_1_10_011_111_100_0_x_00;
      patterns[6034] = 33'b1010110000110111_1_1_10_011_111_100_0_x_00;
      patterns[6035] = 33'b1010110000110111_0_0_00_000_000_000_0_0_00;
      patterns[6036] = 33'b1011010000110111_0_1_11_011_111_100_0_x_00;
      patterns[6037] = 33'b1011110000110111_1_1_11_011_111_100_0_x_00;
      patterns[6038] = 33'b1011110000110111_0_0_00_000_000_000_0_0_00;
      patterns[6039] = 33'b0101010000110000_0_1_xx_011_xxx_100_0_1_01;
      patterns[6040] = 33'b0101110000110000_1_1_xx_011_xxx_100_0_1_01;
      patterns[6041] = 33'b0101110000110000_0_0_00_000_000_000_0_0_00;
      patterns[6042] = 33'b0100010000110000_0_0_xx_011_100_xxx_1_x_xx;
      patterns[6043] = 33'b0100110000110000_1_0_xx_011_100_xxx_1_x_xx;
      patterns[6044] = 33'b0100110000110000_0_0_00_000_000_000_0_0_00;
      patterns[6045] = 33'b0000010001001100_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6046] = 33'b0000110001001100_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6047] = 33'b0000110001001100_0_0_00_000_000_000_0_0_00;
      patterns[6048] = 33'b1000010001000000_0_1_00_100_000_100_0_x_00;
      patterns[6049] = 33'b1000110001000000_1_1_00_100_000_100_0_x_00;
      patterns[6050] = 33'b1000110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6051] = 33'b1001010001000000_0_1_01_100_000_100_0_x_00;
      patterns[6052] = 33'b1001110001000000_1_1_01_100_000_100_0_x_00;
      patterns[6053] = 33'b1001110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6054] = 33'b1010010001000000_0_1_10_100_000_100_0_x_00;
      patterns[6055] = 33'b1010110001000000_1_1_10_100_000_100_0_x_00;
      patterns[6056] = 33'b1010110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6057] = 33'b1011010001000000_0_1_11_100_000_100_0_x_00;
      patterns[6058] = 33'b1011110001000000_1_1_11_100_000_100_0_x_00;
      patterns[6059] = 33'b1011110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6060] = 33'b0101010001000000_0_1_xx_100_xxx_100_0_1_01;
      patterns[6061] = 33'b0101110001000000_1_1_xx_100_xxx_100_0_1_01;
      patterns[6062] = 33'b0101110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6063] = 33'b0100010001000000_0_0_xx_100_100_xxx_1_x_xx;
      patterns[6064] = 33'b0100110001000000_1_0_xx_100_100_xxx_1_x_xx;
      patterns[6065] = 33'b0100110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6066] = 33'b0000010010101000_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6067] = 33'b0000110010101000_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6068] = 33'b0000110010101000_0_0_00_000_000_000_0_0_00;
      patterns[6069] = 33'b1000010001000001_0_1_00_100_001_100_0_x_00;
      patterns[6070] = 33'b1000110001000001_1_1_00_100_001_100_0_x_00;
      patterns[6071] = 33'b1000110001000001_0_0_00_000_000_000_0_0_00;
      patterns[6072] = 33'b1001010001000001_0_1_01_100_001_100_0_x_00;
      patterns[6073] = 33'b1001110001000001_1_1_01_100_001_100_0_x_00;
      patterns[6074] = 33'b1001110001000001_0_0_00_000_000_000_0_0_00;
      patterns[6075] = 33'b1010010001000001_0_1_10_100_001_100_0_x_00;
      patterns[6076] = 33'b1010110001000001_1_1_10_100_001_100_0_x_00;
      patterns[6077] = 33'b1010110001000001_0_0_00_000_000_000_0_0_00;
      patterns[6078] = 33'b1011010001000001_0_1_11_100_001_100_0_x_00;
      patterns[6079] = 33'b1011110001000001_1_1_11_100_001_100_0_x_00;
      patterns[6080] = 33'b1011110001000001_0_0_00_000_000_000_0_0_00;
      patterns[6081] = 33'b0101010001000000_0_1_xx_100_xxx_100_0_1_01;
      patterns[6082] = 33'b0101110001000000_1_1_xx_100_xxx_100_0_1_01;
      patterns[6083] = 33'b0101110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6084] = 33'b0100010001000000_0_0_xx_100_100_xxx_1_x_xx;
      patterns[6085] = 33'b0100110001000000_1_0_xx_100_100_xxx_1_x_xx;
      patterns[6086] = 33'b0100110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6087] = 33'b0000010001000100_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6088] = 33'b0000110001000100_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6089] = 33'b0000110001000100_0_0_00_000_000_000_0_0_00;
      patterns[6090] = 33'b1000010001000010_0_1_00_100_010_100_0_x_00;
      patterns[6091] = 33'b1000110001000010_1_1_00_100_010_100_0_x_00;
      patterns[6092] = 33'b1000110001000010_0_0_00_000_000_000_0_0_00;
      patterns[6093] = 33'b1001010001000010_0_1_01_100_010_100_0_x_00;
      patterns[6094] = 33'b1001110001000010_1_1_01_100_010_100_0_x_00;
      patterns[6095] = 33'b1001110001000010_0_0_00_000_000_000_0_0_00;
      patterns[6096] = 33'b1010010001000010_0_1_10_100_010_100_0_x_00;
      patterns[6097] = 33'b1010110001000010_1_1_10_100_010_100_0_x_00;
      patterns[6098] = 33'b1010110001000010_0_0_00_000_000_000_0_0_00;
      patterns[6099] = 33'b1011010001000010_0_1_11_100_010_100_0_x_00;
      patterns[6100] = 33'b1011110001000010_1_1_11_100_010_100_0_x_00;
      patterns[6101] = 33'b1011110001000010_0_0_00_000_000_000_0_0_00;
      patterns[6102] = 33'b0101010001000000_0_1_xx_100_xxx_100_0_1_01;
      patterns[6103] = 33'b0101110001000000_1_1_xx_100_xxx_100_0_1_01;
      patterns[6104] = 33'b0101110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6105] = 33'b0100010001000000_0_0_xx_100_100_xxx_1_x_xx;
      patterns[6106] = 33'b0100110001000000_1_0_xx_100_100_xxx_1_x_xx;
      patterns[6107] = 33'b0100110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6108] = 33'b0000010000111001_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6109] = 33'b0000110000111001_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6110] = 33'b0000110000111001_0_0_00_000_000_000_0_0_00;
      patterns[6111] = 33'b1000010001000011_0_1_00_100_011_100_0_x_00;
      patterns[6112] = 33'b1000110001000011_1_1_00_100_011_100_0_x_00;
      patterns[6113] = 33'b1000110001000011_0_0_00_000_000_000_0_0_00;
      patterns[6114] = 33'b1001010001000011_0_1_01_100_011_100_0_x_00;
      patterns[6115] = 33'b1001110001000011_1_1_01_100_011_100_0_x_00;
      patterns[6116] = 33'b1001110001000011_0_0_00_000_000_000_0_0_00;
      patterns[6117] = 33'b1010010001000011_0_1_10_100_011_100_0_x_00;
      patterns[6118] = 33'b1010110001000011_1_1_10_100_011_100_0_x_00;
      patterns[6119] = 33'b1010110001000011_0_0_00_000_000_000_0_0_00;
      patterns[6120] = 33'b1011010001000011_0_1_11_100_011_100_0_x_00;
      patterns[6121] = 33'b1011110001000011_1_1_11_100_011_100_0_x_00;
      patterns[6122] = 33'b1011110001000011_0_0_00_000_000_000_0_0_00;
      patterns[6123] = 33'b0101010001000000_0_1_xx_100_xxx_100_0_1_01;
      patterns[6124] = 33'b0101110001000000_1_1_xx_100_xxx_100_0_1_01;
      patterns[6125] = 33'b0101110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6126] = 33'b0100010001000000_0_0_xx_100_100_xxx_1_x_xx;
      patterns[6127] = 33'b0100110001000000_1_0_xx_100_100_xxx_1_x_xx;
      patterns[6128] = 33'b0100110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6129] = 33'b0000010000010010_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6130] = 33'b0000110000010010_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6131] = 33'b0000110000010010_0_0_00_000_000_000_0_0_00;
      patterns[6132] = 33'b1000010001000100_0_1_00_100_100_100_0_x_00;
      patterns[6133] = 33'b1000110001000100_1_1_00_100_100_100_0_x_00;
      patterns[6134] = 33'b1000110001000100_0_0_00_000_000_000_0_0_00;
      patterns[6135] = 33'b1001010001000100_0_1_01_100_100_100_0_x_00;
      patterns[6136] = 33'b1001110001000100_1_1_01_100_100_100_0_x_00;
      patterns[6137] = 33'b1001110001000100_0_0_00_000_000_000_0_0_00;
      patterns[6138] = 33'b1010010001000100_0_1_10_100_100_100_0_x_00;
      patterns[6139] = 33'b1010110001000100_1_1_10_100_100_100_0_x_00;
      patterns[6140] = 33'b1010110001000100_0_0_00_000_000_000_0_0_00;
      patterns[6141] = 33'b1011010001000100_0_1_11_100_100_100_0_x_00;
      patterns[6142] = 33'b1011110001000100_1_1_11_100_100_100_0_x_00;
      patterns[6143] = 33'b1011110001000100_0_0_00_000_000_000_0_0_00;
      patterns[6144] = 33'b0101010001000000_0_1_xx_100_xxx_100_0_1_01;
      patterns[6145] = 33'b0101110001000000_1_1_xx_100_xxx_100_0_1_01;
      patterns[6146] = 33'b0101110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6147] = 33'b0100010001000000_0_0_xx_100_100_xxx_1_x_xx;
      patterns[6148] = 33'b0100110001000000_1_0_xx_100_100_xxx_1_x_xx;
      patterns[6149] = 33'b0100110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6150] = 33'b0000010000011000_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6151] = 33'b0000110000011000_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6152] = 33'b0000110000011000_0_0_00_000_000_000_0_0_00;
      patterns[6153] = 33'b1000010001000101_0_1_00_100_101_100_0_x_00;
      patterns[6154] = 33'b1000110001000101_1_1_00_100_101_100_0_x_00;
      patterns[6155] = 33'b1000110001000101_0_0_00_000_000_000_0_0_00;
      patterns[6156] = 33'b1001010001000101_0_1_01_100_101_100_0_x_00;
      patterns[6157] = 33'b1001110001000101_1_1_01_100_101_100_0_x_00;
      patterns[6158] = 33'b1001110001000101_0_0_00_000_000_000_0_0_00;
      patterns[6159] = 33'b1010010001000101_0_1_10_100_101_100_0_x_00;
      patterns[6160] = 33'b1010110001000101_1_1_10_100_101_100_0_x_00;
      patterns[6161] = 33'b1010110001000101_0_0_00_000_000_000_0_0_00;
      patterns[6162] = 33'b1011010001000101_0_1_11_100_101_100_0_x_00;
      patterns[6163] = 33'b1011110001000101_1_1_11_100_101_100_0_x_00;
      patterns[6164] = 33'b1011110001000101_0_0_00_000_000_000_0_0_00;
      patterns[6165] = 33'b0101010001000000_0_1_xx_100_xxx_100_0_1_01;
      patterns[6166] = 33'b0101110001000000_1_1_xx_100_xxx_100_0_1_01;
      patterns[6167] = 33'b0101110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6168] = 33'b0100010001000000_0_0_xx_100_100_xxx_1_x_xx;
      patterns[6169] = 33'b0100110001000000_1_0_xx_100_100_xxx_1_x_xx;
      patterns[6170] = 33'b0100110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6171] = 33'b0000010000111001_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6172] = 33'b0000110000111001_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6173] = 33'b0000110000111001_0_0_00_000_000_000_0_0_00;
      patterns[6174] = 33'b1000010001000110_0_1_00_100_110_100_0_x_00;
      patterns[6175] = 33'b1000110001000110_1_1_00_100_110_100_0_x_00;
      patterns[6176] = 33'b1000110001000110_0_0_00_000_000_000_0_0_00;
      patterns[6177] = 33'b1001010001000110_0_1_01_100_110_100_0_x_00;
      patterns[6178] = 33'b1001110001000110_1_1_01_100_110_100_0_x_00;
      patterns[6179] = 33'b1001110001000110_0_0_00_000_000_000_0_0_00;
      patterns[6180] = 33'b1010010001000110_0_1_10_100_110_100_0_x_00;
      patterns[6181] = 33'b1010110001000110_1_1_10_100_110_100_0_x_00;
      patterns[6182] = 33'b1010110001000110_0_0_00_000_000_000_0_0_00;
      patterns[6183] = 33'b1011010001000110_0_1_11_100_110_100_0_x_00;
      patterns[6184] = 33'b1011110001000110_1_1_11_100_110_100_0_x_00;
      patterns[6185] = 33'b1011110001000110_0_0_00_000_000_000_0_0_00;
      patterns[6186] = 33'b0101010001000000_0_1_xx_100_xxx_100_0_1_01;
      patterns[6187] = 33'b0101110001000000_1_1_xx_100_xxx_100_0_1_01;
      patterns[6188] = 33'b0101110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6189] = 33'b0100010001000000_0_0_xx_100_100_xxx_1_x_xx;
      patterns[6190] = 33'b0100110001000000_1_0_xx_100_100_xxx_1_x_xx;
      patterns[6191] = 33'b0100110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6192] = 33'b0000010010101010_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6193] = 33'b0000110010101010_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6194] = 33'b0000110010101010_0_0_00_000_000_000_0_0_00;
      patterns[6195] = 33'b1000010001000111_0_1_00_100_111_100_0_x_00;
      patterns[6196] = 33'b1000110001000111_1_1_00_100_111_100_0_x_00;
      patterns[6197] = 33'b1000110001000111_0_0_00_000_000_000_0_0_00;
      patterns[6198] = 33'b1001010001000111_0_1_01_100_111_100_0_x_00;
      patterns[6199] = 33'b1001110001000111_1_1_01_100_111_100_0_x_00;
      patterns[6200] = 33'b1001110001000111_0_0_00_000_000_000_0_0_00;
      patterns[6201] = 33'b1010010001000111_0_1_10_100_111_100_0_x_00;
      patterns[6202] = 33'b1010110001000111_1_1_10_100_111_100_0_x_00;
      patterns[6203] = 33'b1010110001000111_0_0_00_000_000_000_0_0_00;
      patterns[6204] = 33'b1011010001000111_0_1_11_100_111_100_0_x_00;
      patterns[6205] = 33'b1011110001000111_1_1_11_100_111_100_0_x_00;
      patterns[6206] = 33'b1011110001000111_0_0_00_000_000_000_0_0_00;
      patterns[6207] = 33'b0101010001000000_0_1_xx_100_xxx_100_0_1_01;
      patterns[6208] = 33'b0101110001000000_1_1_xx_100_xxx_100_0_1_01;
      patterns[6209] = 33'b0101110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6210] = 33'b0100010001000000_0_0_xx_100_100_xxx_1_x_xx;
      patterns[6211] = 33'b0100110001000000_1_0_xx_100_100_xxx_1_x_xx;
      patterns[6212] = 33'b0100110001000000_0_0_00_000_000_000_0_0_00;
      patterns[6213] = 33'b0000010000100101_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6214] = 33'b0000110000100101_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6215] = 33'b0000110000100101_0_0_00_000_000_000_0_0_00;
      patterns[6216] = 33'b1000010001010000_0_1_00_101_000_100_0_x_00;
      patterns[6217] = 33'b1000110001010000_1_1_00_101_000_100_0_x_00;
      patterns[6218] = 33'b1000110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6219] = 33'b1001010001010000_0_1_01_101_000_100_0_x_00;
      patterns[6220] = 33'b1001110001010000_1_1_01_101_000_100_0_x_00;
      patterns[6221] = 33'b1001110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6222] = 33'b1010010001010000_0_1_10_101_000_100_0_x_00;
      patterns[6223] = 33'b1010110001010000_1_1_10_101_000_100_0_x_00;
      patterns[6224] = 33'b1010110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6225] = 33'b1011010001010000_0_1_11_101_000_100_0_x_00;
      patterns[6226] = 33'b1011110001010000_1_1_11_101_000_100_0_x_00;
      patterns[6227] = 33'b1011110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6228] = 33'b0101010001010000_0_1_xx_101_xxx_100_0_1_01;
      patterns[6229] = 33'b0101110001010000_1_1_xx_101_xxx_100_0_1_01;
      patterns[6230] = 33'b0101110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6231] = 33'b0100010001010000_0_0_xx_101_100_xxx_1_x_xx;
      patterns[6232] = 33'b0100110001010000_1_0_xx_101_100_xxx_1_x_xx;
      patterns[6233] = 33'b0100110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6234] = 33'b0000010001110100_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6235] = 33'b0000110001110100_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6236] = 33'b0000110001110100_0_0_00_000_000_000_0_0_00;
      patterns[6237] = 33'b1000010001010001_0_1_00_101_001_100_0_x_00;
      patterns[6238] = 33'b1000110001010001_1_1_00_101_001_100_0_x_00;
      patterns[6239] = 33'b1000110001010001_0_0_00_000_000_000_0_0_00;
      patterns[6240] = 33'b1001010001010001_0_1_01_101_001_100_0_x_00;
      patterns[6241] = 33'b1001110001010001_1_1_01_101_001_100_0_x_00;
      patterns[6242] = 33'b1001110001010001_0_0_00_000_000_000_0_0_00;
      patterns[6243] = 33'b1010010001010001_0_1_10_101_001_100_0_x_00;
      patterns[6244] = 33'b1010110001010001_1_1_10_101_001_100_0_x_00;
      patterns[6245] = 33'b1010110001010001_0_0_00_000_000_000_0_0_00;
      patterns[6246] = 33'b1011010001010001_0_1_11_101_001_100_0_x_00;
      patterns[6247] = 33'b1011110001010001_1_1_11_101_001_100_0_x_00;
      patterns[6248] = 33'b1011110001010001_0_0_00_000_000_000_0_0_00;
      patterns[6249] = 33'b0101010001010000_0_1_xx_101_xxx_100_0_1_01;
      patterns[6250] = 33'b0101110001010000_1_1_xx_101_xxx_100_0_1_01;
      patterns[6251] = 33'b0101110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6252] = 33'b0100010001010000_0_0_xx_101_100_xxx_1_x_xx;
      patterns[6253] = 33'b0100110001010000_1_0_xx_101_100_xxx_1_x_xx;
      patterns[6254] = 33'b0100110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6255] = 33'b0000010001100111_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6256] = 33'b0000110001100111_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6257] = 33'b0000110001100111_0_0_00_000_000_000_0_0_00;
      patterns[6258] = 33'b1000010001010010_0_1_00_101_010_100_0_x_00;
      patterns[6259] = 33'b1000110001010010_1_1_00_101_010_100_0_x_00;
      patterns[6260] = 33'b1000110001010010_0_0_00_000_000_000_0_0_00;
      patterns[6261] = 33'b1001010001010010_0_1_01_101_010_100_0_x_00;
      patterns[6262] = 33'b1001110001010010_1_1_01_101_010_100_0_x_00;
      patterns[6263] = 33'b1001110001010010_0_0_00_000_000_000_0_0_00;
      patterns[6264] = 33'b1010010001010010_0_1_10_101_010_100_0_x_00;
      patterns[6265] = 33'b1010110001010010_1_1_10_101_010_100_0_x_00;
      patterns[6266] = 33'b1010110001010010_0_0_00_000_000_000_0_0_00;
      patterns[6267] = 33'b1011010001010010_0_1_11_101_010_100_0_x_00;
      patterns[6268] = 33'b1011110001010010_1_1_11_101_010_100_0_x_00;
      patterns[6269] = 33'b1011110001010010_0_0_00_000_000_000_0_0_00;
      patterns[6270] = 33'b0101010001010000_0_1_xx_101_xxx_100_0_1_01;
      patterns[6271] = 33'b0101110001010000_1_1_xx_101_xxx_100_0_1_01;
      patterns[6272] = 33'b0101110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6273] = 33'b0100010001010000_0_0_xx_101_100_xxx_1_x_xx;
      patterns[6274] = 33'b0100110001010000_1_0_xx_101_100_xxx_1_x_xx;
      patterns[6275] = 33'b0100110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6276] = 33'b0000010001110110_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6277] = 33'b0000110001110110_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6278] = 33'b0000110001110110_0_0_00_000_000_000_0_0_00;
      patterns[6279] = 33'b1000010001010011_0_1_00_101_011_100_0_x_00;
      patterns[6280] = 33'b1000110001010011_1_1_00_101_011_100_0_x_00;
      patterns[6281] = 33'b1000110001010011_0_0_00_000_000_000_0_0_00;
      patterns[6282] = 33'b1001010001010011_0_1_01_101_011_100_0_x_00;
      patterns[6283] = 33'b1001110001010011_1_1_01_101_011_100_0_x_00;
      patterns[6284] = 33'b1001110001010011_0_0_00_000_000_000_0_0_00;
      patterns[6285] = 33'b1010010001010011_0_1_10_101_011_100_0_x_00;
      patterns[6286] = 33'b1010110001010011_1_1_10_101_011_100_0_x_00;
      patterns[6287] = 33'b1010110001010011_0_0_00_000_000_000_0_0_00;
      patterns[6288] = 33'b1011010001010011_0_1_11_101_011_100_0_x_00;
      patterns[6289] = 33'b1011110001010011_1_1_11_101_011_100_0_x_00;
      patterns[6290] = 33'b1011110001010011_0_0_00_000_000_000_0_0_00;
      patterns[6291] = 33'b0101010001010000_0_1_xx_101_xxx_100_0_1_01;
      patterns[6292] = 33'b0101110001010000_1_1_xx_101_xxx_100_0_1_01;
      patterns[6293] = 33'b0101110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6294] = 33'b0100010001010000_0_0_xx_101_100_xxx_1_x_xx;
      patterns[6295] = 33'b0100110001010000_1_0_xx_101_100_xxx_1_x_xx;
      patterns[6296] = 33'b0100110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6297] = 33'b0000010010110110_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6298] = 33'b0000110010110110_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6299] = 33'b0000110010110110_0_0_00_000_000_000_0_0_00;
      patterns[6300] = 33'b1000010001010100_0_1_00_101_100_100_0_x_00;
      patterns[6301] = 33'b1000110001010100_1_1_00_101_100_100_0_x_00;
      patterns[6302] = 33'b1000110001010100_0_0_00_000_000_000_0_0_00;
      patterns[6303] = 33'b1001010001010100_0_1_01_101_100_100_0_x_00;
      patterns[6304] = 33'b1001110001010100_1_1_01_101_100_100_0_x_00;
      patterns[6305] = 33'b1001110001010100_0_0_00_000_000_000_0_0_00;
      patterns[6306] = 33'b1010010001010100_0_1_10_101_100_100_0_x_00;
      patterns[6307] = 33'b1010110001010100_1_1_10_101_100_100_0_x_00;
      patterns[6308] = 33'b1010110001010100_0_0_00_000_000_000_0_0_00;
      patterns[6309] = 33'b1011010001010100_0_1_11_101_100_100_0_x_00;
      patterns[6310] = 33'b1011110001010100_1_1_11_101_100_100_0_x_00;
      patterns[6311] = 33'b1011110001010100_0_0_00_000_000_000_0_0_00;
      patterns[6312] = 33'b0101010001010000_0_1_xx_101_xxx_100_0_1_01;
      patterns[6313] = 33'b0101110001010000_1_1_xx_101_xxx_100_0_1_01;
      patterns[6314] = 33'b0101110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6315] = 33'b0100010001010000_0_0_xx_101_100_xxx_1_x_xx;
      patterns[6316] = 33'b0100110001010000_1_0_xx_101_100_xxx_1_x_xx;
      patterns[6317] = 33'b0100110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6318] = 33'b0000010010101100_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6319] = 33'b0000110010101100_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6320] = 33'b0000110010101100_0_0_00_000_000_000_0_0_00;
      patterns[6321] = 33'b1000010001010101_0_1_00_101_101_100_0_x_00;
      patterns[6322] = 33'b1000110001010101_1_1_00_101_101_100_0_x_00;
      patterns[6323] = 33'b1000110001010101_0_0_00_000_000_000_0_0_00;
      patterns[6324] = 33'b1001010001010101_0_1_01_101_101_100_0_x_00;
      patterns[6325] = 33'b1001110001010101_1_1_01_101_101_100_0_x_00;
      patterns[6326] = 33'b1001110001010101_0_0_00_000_000_000_0_0_00;
      patterns[6327] = 33'b1010010001010101_0_1_10_101_101_100_0_x_00;
      patterns[6328] = 33'b1010110001010101_1_1_10_101_101_100_0_x_00;
      patterns[6329] = 33'b1010110001010101_0_0_00_000_000_000_0_0_00;
      patterns[6330] = 33'b1011010001010101_0_1_11_101_101_100_0_x_00;
      patterns[6331] = 33'b1011110001010101_1_1_11_101_101_100_0_x_00;
      patterns[6332] = 33'b1011110001010101_0_0_00_000_000_000_0_0_00;
      patterns[6333] = 33'b0101010001010000_0_1_xx_101_xxx_100_0_1_01;
      patterns[6334] = 33'b0101110001010000_1_1_xx_101_xxx_100_0_1_01;
      patterns[6335] = 33'b0101110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6336] = 33'b0100010001010000_0_0_xx_101_100_xxx_1_x_xx;
      patterns[6337] = 33'b0100110001010000_1_0_xx_101_100_xxx_1_x_xx;
      patterns[6338] = 33'b0100110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6339] = 33'b0000010010001101_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6340] = 33'b0000110010001101_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6341] = 33'b0000110010001101_0_0_00_000_000_000_0_0_00;
      patterns[6342] = 33'b1000010001010110_0_1_00_101_110_100_0_x_00;
      patterns[6343] = 33'b1000110001010110_1_1_00_101_110_100_0_x_00;
      patterns[6344] = 33'b1000110001010110_0_0_00_000_000_000_0_0_00;
      patterns[6345] = 33'b1001010001010110_0_1_01_101_110_100_0_x_00;
      patterns[6346] = 33'b1001110001010110_1_1_01_101_110_100_0_x_00;
      patterns[6347] = 33'b1001110001010110_0_0_00_000_000_000_0_0_00;
      patterns[6348] = 33'b1010010001010110_0_1_10_101_110_100_0_x_00;
      patterns[6349] = 33'b1010110001010110_1_1_10_101_110_100_0_x_00;
      patterns[6350] = 33'b1010110001010110_0_0_00_000_000_000_0_0_00;
      patterns[6351] = 33'b1011010001010110_0_1_11_101_110_100_0_x_00;
      patterns[6352] = 33'b1011110001010110_1_1_11_101_110_100_0_x_00;
      patterns[6353] = 33'b1011110001010110_0_0_00_000_000_000_0_0_00;
      patterns[6354] = 33'b0101010001010000_0_1_xx_101_xxx_100_0_1_01;
      patterns[6355] = 33'b0101110001010000_1_1_xx_101_xxx_100_0_1_01;
      patterns[6356] = 33'b0101110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6357] = 33'b0100010001010000_0_0_xx_101_100_xxx_1_x_xx;
      patterns[6358] = 33'b0100110001010000_1_0_xx_101_100_xxx_1_x_xx;
      patterns[6359] = 33'b0100110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6360] = 33'b0000010011111110_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6361] = 33'b0000110011111110_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6362] = 33'b0000110011111110_0_0_00_000_000_000_0_0_00;
      patterns[6363] = 33'b1000010001010111_0_1_00_101_111_100_0_x_00;
      patterns[6364] = 33'b1000110001010111_1_1_00_101_111_100_0_x_00;
      patterns[6365] = 33'b1000110001010111_0_0_00_000_000_000_0_0_00;
      patterns[6366] = 33'b1001010001010111_0_1_01_101_111_100_0_x_00;
      patterns[6367] = 33'b1001110001010111_1_1_01_101_111_100_0_x_00;
      patterns[6368] = 33'b1001110001010111_0_0_00_000_000_000_0_0_00;
      patterns[6369] = 33'b1010010001010111_0_1_10_101_111_100_0_x_00;
      patterns[6370] = 33'b1010110001010111_1_1_10_101_111_100_0_x_00;
      patterns[6371] = 33'b1010110001010111_0_0_00_000_000_000_0_0_00;
      patterns[6372] = 33'b1011010001010111_0_1_11_101_111_100_0_x_00;
      patterns[6373] = 33'b1011110001010111_1_1_11_101_111_100_0_x_00;
      patterns[6374] = 33'b1011110001010111_0_0_00_000_000_000_0_0_00;
      patterns[6375] = 33'b0101010001010000_0_1_xx_101_xxx_100_0_1_01;
      patterns[6376] = 33'b0101110001010000_1_1_xx_101_xxx_100_0_1_01;
      patterns[6377] = 33'b0101110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6378] = 33'b0100010001010000_0_0_xx_101_100_xxx_1_x_xx;
      patterns[6379] = 33'b0100110001010000_1_0_xx_101_100_xxx_1_x_xx;
      patterns[6380] = 33'b0100110001010000_0_0_00_000_000_000_0_0_00;
      patterns[6381] = 33'b0000010001011110_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6382] = 33'b0000110001011110_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6383] = 33'b0000110001011110_0_0_00_000_000_000_0_0_00;
      patterns[6384] = 33'b1000010001100000_0_1_00_110_000_100_0_x_00;
      patterns[6385] = 33'b1000110001100000_1_1_00_110_000_100_0_x_00;
      patterns[6386] = 33'b1000110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6387] = 33'b1001010001100000_0_1_01_110_000_100_0_x_00;
      patterns[6388] = 33'b1001110001100000_1_1_01_110_000_100_0_x_00;
      patterns[6389] = 33'b1001110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6390] = 33'b1010010001100000_0_1_10_110_000_100_0_x_00;
      patterns[6391] = 33'b1010110001100000_1_1_10_110_000_100_0_x_00;
      patterns[6392] = 33'b1010110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6393] = 33'b1011010001100000_0_1_11_110_000_100_0_x_00;
      patterns[6394] = 33'b1011110001100000_1_1_11_110_000_100_0_x_00;
      patterns[6395] = 33'b1011110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6396] = 33'b0101010001100000_0_1_xx_110_xxx_100_0_1_01;
      patterns[6397] = 33'b0101110001100000_1_1_xx_110_xxx_100_0_1_01;
      patterns[6398] = 33'b0101110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6399] = 33'b0100010001100000_0_0_xx_110_100_xxx_1_x_xx;
      patterns[6400] = 33'b0100110001100000_1_0_xx_110_100_xxx_1_x_xx;
      patterns[6401] = 33'b0100110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6402] = 33'b0000010001100110_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6403] = 33'b0000110001100110_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6404] = 33'b0000110001100110_0_0_00_000_000_000_0_0_00;
      patterns[6405] = 33'b1000010001100001_0_1_00_110_001_100_0_x_00;
      patterns[6406] = 33'b1000110001100001_1_1_00_110_001_100_0_x_00;
      patterns[6407] = 33'b1000110001100001_0_0_00_000_000_000_0_0_00;
      patterns[6408] = 33'b1001010001100001_0_1_01_110_001_100_0_x_00;
      patterns[6409] = 33'b1001110001100001_1_1_01_110_001_100_0_x_00;
      patterns[6410] = 33'b1001110001100001_0_0_00_000_000_000_0_0_00;
      patterns[6411] = 33'b1010010001100001_0_1_10_110_001_100_0_x_00;
      patterns[6412] = 33'b1010110001100001_1_1_10_110_001_100_0_x_00;
      patterns[6413] = 33'b1010110001100001_0_0_00_000_000_000_0_0_00;
      patterns[6414] = 33'b1011010001100001_0_1_11_110_001_100_0_x_00;
      patterns[6415] = 33'b1011110001100001_1_1_11_110_001_100_0_x_00;
      patterns[6416] = 33'b1011110001100001_0_0_00_000_000_000_0_0_00;
      patterns[6417] = 33'b0101010001100000_0_1_xx_110_xxx_100_0_1_01;
      patterns[6418] = 33'b0101110001100000_1_1_xx_110_xxx_100_0_1_01;
      patterns[6419] = 33'b0101110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6420] = 33'b0100010001100000_0_0_xx_110_100_xxx_1_x_xx;
      patterns[6421] = 33'b0100110001100000_1_0_xx_110_100_xxx_1_x_xx;
      patterns[6422] = 33'b0100110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6423] = 33'b0000010011100110_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6424] = 33'b0000110011100110_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6425] = 33'b0000110011100110_0_0_00_000_000_000_0_0_00;
      patterns[6426] = 33'b1000010001100010_0_1_00_110_010_100_0_x_00;
      patterns[6427] = 33'b1000110001100010_1_1_00_110_010_100_0_x_00;
      patterns[6428] = 33'b1000110001100010_0_0_00_000_000_000_0_0_00;
      patterns[6429] = 33'b1001010001100010_0_1_01_110_010_100_0_x_00;
      patterns[6430] = 33'b1001110001100010_1_1_01_110_010_100_0_x_00;
      patterns[6431] = 33'b1001110001100010_0_0_00_000_000_000_0_0_00;
      patterns[6432] = 33'b1010010001100010_0_1_10_110_010_100_0_x_00;
      patterns[6433] = 33'b1010110001100010_1_1_10_110_010_100_0_x_00;
      patterns[6434] = 33'b1010110001100010_0_0_00_000_000_000_0_0_00;
      patterns[6435] = 33'b1011010001100010_0_1_11_110_010_100_0_x_00;
      patterns[6436] = 33'b1011110001100010_1_1_11_110_010_100_0_x_00;
      patterns[6437] = 33'b1011110001100010_0_0_00_000_000_000_0_0_00;
      patterns[6438] = 33'b0101010001100000_0_1_xx_110_xxx_100_0_1_01;
      patterns[6439] = 33'b0101110001100000_1_1_xx_110_xxx_100_0_1_01;
      patterns[6440] = 33'b0101110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6441] = 33'b0100010001100000_0_0_xx_110_100_xxx_1_x_xx;
      patterns[6442] = 33'b0100110001100000_1_0_xx_110_100_xxx_1_x_xx;
      patterns[6443] = 33'b0100110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6444] = 33'b0000010010101001_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6445] = 33'b0000110010101001_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6446] = 33'b0000110010101001_0_0_00_000_000_000_0_0_00;
      patterns[6447] = 33'b1000010001100011_0_1_00_110_011_100_0_x_00;
      patterns[6448] = 33'b1000110001100011_1_1_00_110_011_100_0_x_00;
      patterns[6449] = 33'b1000110001100011_0_0_00_000_000_000_0_0_00;
      patterns[6450] = 33'b1001010001100011_0_1_01_110_011_100_0_x_00;
      patterns[6451] = 33'b1001110001100011_1_1_01_110_011_100_0_x_00;
      patterns[6452] = 33'b1001110001100011_0_0_00_000_000_000_0_0_00;
      patterns[6453] = 33'b1010010001100011_0_1_10_110_011_100_0_x_00;
      patterns[6454] = 33'b1010110001100011_1_1_10_110_011_100_0_x_00;
      patterns[6455] = 33'b1010110001100011_0_0_00_000_000_000_0_0_00;
      patterns[6456] = 33'b1011010001100011_0_1_11_110_011_100_0_x_00;
      patterns[6457] = 33'b1011110001100011_1_1_11_110_011_100_0_x_00;
      patterns[6458] = 33'b1011110001100011_0_0_00_000_000_000_0_0_00;
      patterns[6459] = 33'b0101010001100000_0_1_xx_110_xxx_100_0_1_01;
      patterns[6460] = 33'b0101110001100000_1_1_xx_110_xxx_100_0_1_01;
      patterns[6461] = 33'b0101110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6462] = 33'b0100010001100000_0_0_xx_110_100_xxx_1_x_xx;
      patterns[6463] = 33'b0100110001100000_1_0_xx_110_100_xxx_1_x_xx;
      patterns[6464] = 33'b0100110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6465] = 33'b0000010010101011_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6466] = 33'b0000110010101011_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6467] = 33'b0000110010101011_0_0_00_000_000_000_0_0_00;
      patterns[6468] = 33'b1000010001100100_0_1_00_110_100_100_0_x_00;
      patterns[6469] = 33'b1000110001100100_1_1_00_110_100_100_0_x_00;
      patterns[6470] = 33'b1000110001100100_0_0_00_000_000_000_0_0_00;
      patterns[6471] = 33'b1001010001100100_0_1_01_110_100_100_0_x_00;
      patterns[6472] = 33'b1001110001100100_1_1_01_110_100_100_0_x_00;
      patterns[6473] = 33'b1001110001100100_0_0_00_000_000_000_0_0_00;
      patterns[6474] = 33'b1010010001100100_0_1_10_110_100_100_0_x_00;
      patterns[6475] = 33'b1010110001100100_1_1_10_110_100_100_0_x_00;
      patterns[6476] = 33'b1010110001100100_0_0_00_000_000_000_0_0_00;
      patterns[6477] = 33'b1011010001100100_0_1_11_110_100_100_0_x_00;
      patterns[6478] = 33'b1011110001100100_1_1_11_110_100_100_0_x_00;
      patterns[6479] = 33'b1011110001100100_0_0_00_000_000_000_0_0_00;
      patterns[6480] = 33'b0101010001100000_0_1_xx_110_xxx_100_0_1_01;
      patterns[6481] = 33'b0101110001100000_1_1_xx_110_xxx_100_0_1_01;
      patterns[6482] = 33'b0101110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6483] = 33'b0100010001100000_0_0_xx_110_100_xxx_1_x_xx;
      patterns[6484] = 33'b0100110001100000_1_0_xx_110_100_xxx_1_x_xx;
      patterns[6485] = 33'b0100110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6486] = 33'b0000010011101111_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6487] = 33'b0000110011101111_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6488] = 33'b0000110011101111_0_0_00_000_000_000_0_0_00;
      patterns[6489] = 33'b1000010001100101_0_1_00_110_101_100_0_x_00;
      patterns[6490] = 33'b1000110001100101_1_1_00_110_101_100_0_x_00;
      patterns[6491] = 33'b1000110001100101_0_0_00_000_000_000_0_0_00;
      patterns[6492] = 33'b1001010001100101_0_1_01_110_101_100_0_x_00;
      patterns[6493] = 33'b1001110001100101_1_1_01_110_101_100_0_x_00;
      patterns[6494] = 33'b1001110001100101_0_0_00_000_000_000_0_0_00;
      patterns[6495] = 33'b1010010001100101_0_1_10_110_101_100_0_x_00;
      patterns[6496] = 33'b1010110001100101_1_1_10_110_101_100_0_x_00;
      patterns[6497] = 33'b1010110001100101_0_0_00_000_000_000_0_0_00;
      patterns[6498] = 33'b1011010001100101_0_1_11_110_101_100_0_x_00;
      patterns[6499] = 33'b1011110001100101_1_1_11_110_101_100_0_x_00;
      patterns[6500] = 33'b1011110001100101_0_0_00_000_000_000_0_0_00;
      patterns[6501] = 33'b0101010001100000_0_1_xx_110_xxx_100_0_1_01;
      patterns[6502] = 33'b0101110001100000_1_1_xx_110_xxx_100_0_1_01;
      patterns[6503] = 33'b0101110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6504] = 33'b0100010001100000_0_0_xx_110_100_xxx_1_x_xx;
      patterns[6505] = 33'b0100110001100000_1_0_xx_110_100_xxx_1_x_xx;
      patterns[6506] = 33'b0100110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6507] = 33'b0000010001110100_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6508] = 33'b0000110001110100_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6509] = 33'b0000110001110100_0_0_00_000_000_000_0_0_00;
      patterns[6510] = 33'b1000010001100110_0_1_00_110_110_100_0_x_00;
      patterns[6511] = 33'b1000110001100110_1_1_00_110_110_100_0_x_00;
      patterns[6512] = 33'b1000110001100110_0_0_00_000_000_000_0_0_00;
      patterns[6513] = 33'b1001010001100110_0_1_01_110_110_100_0_x_00;
      patterns[6514] = 33'b1001110001100110_1_1_01_110_110_100_0_x_00;
      patterns[6515] = 33'b1001110001100110_0_0_00_000_000_000_0_0_00;
      patterns[6516] = 33'b1010010001100110_0_1_10_110_110_100_0_x_00;
      patterns[6517] = 33'b1010110001100110_1_1_10_110_110_100_0_x_00;
      patterns[6518] = 33'b1010110001100110_0_0_00_000_000_000_0_0_00;
      patterns[6519] = 33'b1011010001100110_0_1_11_110_110_100_0_x_00;
      patterns[6520] = 33'b1011110001100110_1_1_11_110_110_100_0_x_00;
      patterns[6521] = 33'b1011110001100110_0_0_00_000_000_000_0_0_00;
      patterns[6522] = 33'b0101010001100000_0_1_xx_110_xxx_100_0_1_01;
      patterns[6523] = 33'b0101110001100000_1_1_xx_110_xxx_100_0_1_01;
      patterns[6524] = 33'b0101110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6525] = 33'b0100010001100000_0_0_xx_110_100_xxx_1_x_xx;
      patterns[6526] = 33'b0100110001100000_1_0_xx_110_100_xxx_1_x_xx;
      patterns[6527] = 33'b0100110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6528] = 33'b0000010011100001_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6529] = 33'b0000110011100001_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6530] = 33'b0000110011100001_0_0_00_000_000_000_0_0_00;
      patterns[6531] = 33'b1000010001100111_0_1_00_110_111_100_0_x_00;
      patterns[6532] = 33'b1000110001100111_1_1_00_110_111_100_0_x_00;
      patterns[6533] = 33'b1000110001100111_0_0_00_000_000_000_0_0_00;
      patterns[6534] = 33'b1001010001100111_0_1_01_110_111_100_0_x_00;
      patterns[6535] = 33'b1001110001100111_1_1_01_110_111_100_0_x_00;
      patterns[6536] = 33'b1001110001100111_0_0_00_000_000_000_0_0_00;
      patterns[6537] = 33'b1010010001100111_0_1_10_110_111_100_0_x_00;
      patterns[6538] = 33'b1010110001100111_1_1_10_110_111_100_0_x_00;
      patterns[6539] = 33'b1010110001100111_0_0_00_000_000_000_0_0_00;
      patterns[6540] = 33'b1011010001100111_0_1_11_110_111_100_0_x_00;
      patterns[6541] = 33'b1011110001100111_1_1_11_110_111_100_0_x_00;
      patterns[6542] = 33'b1011110001100111_0_0_00_000_000_000_0_0_00;
      patterns[6543] = 33'b0101010001100000_0_1_xx_110_xxx_100_0_1_01;
      patterns[6544] = 33'b0101110001100000_1_1_xx_110_xxx_100_0_1_01;
      patterns[6545] = 33'b0101110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6546] = 33'b0100010001100000_0_0_xx_110_100_xxx_1_x_xx;
      patterns[6547] = 33'b0100110001100000_1_0_xx_110_100_xxx_1_x_xx;
      patterns[6548] = 33'b0100110001100000_0_0_00_000_000_000_0_0_00;
      patterns[6549] = 33'b0000010011110011_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6550] = 33'b0000110011110011_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6551] = 33'b0000110011110011_0_0_00_000_000_000_0_0_00;
      patterns[6552] = 33'b1000010001110000_0_1_00_111_000_100_0_x_00;
      patterns[6553] = 33'b1000110001110000_1_1_00_111_000_100_0_x_00;
      patterns[6554] = 33'b1000110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6555] = 33'b1001010001110000_0_1_01_111_000_100_0_x_00;
      patterns[6556] = 33'b1001110001110000_1_1_01_111_000_100_0_x_00;
      patterns[6557] = 33'b1001110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6558] = 33'b1010010001110000_0_1_10_111_000_100_0_x_00;
      patterns[6559] = 33'b1010110001110000_1_1_10_111_000_100_0_x_00;
      patterns[6560] = 33'b1010110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6561] = 33'b1011010001110000_0_1_11_111_000_100_0_x_00;
      patterns[6562] = 33'b1011110001110000_1_1_11_111_000_100_0_x_00;
      patterns[6563] = 33'b1011110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6564] = 33'b0101010001110000_0_1_xx_111_xxx_100_0_1_01;
      patterns[6565] = 33'b0101110001110000_1_1_xx_111_xxx_100_0_1_01;
      patterns[6566] = 33'b0101110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6567] = 33'b0100010001110000_0_0_xx_111_100_xxx_1_x_xx;
      patterns[6568] = 33'b0100110001110000_1_0_xx_111_100_xxx_1_x_xx;
      patterns[6569] = 33'b0100110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6570] = 33'b0000010000001010_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6571] = 33'b0000110000001010_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6572] = 33'b0000110000001010_0_0_00_000_000_000_0_0_00;
      patterns[6573] = 33'b1000010001110001_0_1_00_111_001_100_0_x_00;
      patterns[6574] = 33'b1000110001110001_1_1_00_111_001_100_0_x_00;
      patterns[6575] = 33'b1000110001110001_0_0_00_000_000_000_0_0_00;
      patterns[6576] = 33'b1001010001110001_0_1_01_111_001_100_0_x_00;
      patterns[6577] = 33'b1001110001110001_1_1_01_111_001_100_0_x_00;
      patterns[6578] = 33'b1001110001110001_0_0_00_000_000_000_0_0_00;
      patterns[6579] = 33'b1010010001110001_0_1_10_111_001_100_0_x_00;
      patterns[6580] = 33'b1010110001110001_1_1_10_111_001_100_0_x_00;
      patterns[6581] = 33'b1010110001110001_0_0_00_000_000_000_0_0_00;
      patterns[6582] = 33'b1011010001110001_0_1_11_111_001_100_0_x_00;
      patterns[6583] = 33'b1011110001110001_1_1_11_111_001_100_0_x_00;
      patterns[6584] = 33'b1011110001110001_0_0_00_000_000_000_0_0_00;
      patterns[6585] = 33'b0101010001110000_0_1_xx_111_xxx_100_0_1_01;
      patterns[6586] = 33'b0101110001110000_1_1_xx_111_xxx_100_0_1_01;
      patterns[6587] = 33'b0101110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6588] = 33'b0100010001110000_0_0_xx_111_100_xxx_1_x_xx;
      patterns[6589] = 33'b0100110001110000_1_0_xx_111_100_xxx_1_x_xx;
      patterns[6590] = 33'b0100110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6591] = 33'b0000010011101100_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6592] = 33'b0000110011101100_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6593] = 33'b0000110011101100_0_0_00_000_000_000_0_0_00;
      patterns[6594] = 33'b1000010001110010_0_1_00_111_010_100_0_x_00;
      patterns[6595] = 33'b1000110001110010_1_1_00_111_010_100_0_x_00;
      patterns[6596] = 33'b1000110001110010_0_0_00_000_000_000_0_0_00;
      patterns[6597] = 33'b1001010001110010_0_1_01_111_010_100_0_x_00;
      patterns[6598] = 33'b1001110001110010_1_1_01_111_010_100_0_x_00;
      patterns[6599] = 33'b1001110001110010_0_0_00_000_000_000_0_0_00;
      patterns[6600] = 33'b1010010001110010_0_1_10_111_010_100_0_x_00;
      patterns[6601] = 33'b1010110001110010_1_1_10_111_010_100_0_x_00;
      patterns[6602] = 33'b1010110001110010_0_0_00_000_000_000_0_0_00;
      patterns[6603] = 33'b1011010001110010_0_1_11_111_010_100_0_x_00;
      patterns[6604] = 33'b1011110001110010_1_1_11_111_010_100_0_x_00;
      patterns[6605] = 33'b1011110001110010_0_0_00_000_000_000_0_0_00;
      patterns[6606] = 33'b0101010001110000_0_1_xx_111_xxx_100_0_1_01;
      patterns[6607] = 33'b0101110001110000_1_1_xx_111_xxx_100_0_1_01;
      patterns[6608] = 33'b0101110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6609] = 33'b0100010001110000_0_0_xx_111_100_xxx_1_x_xx;
      patterns[6610] = 33'b0100110001110000_1_0_xx_111_100_xxx_1_x_xx;
      patterns[6611] = 33'b0100110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6612] = 33'b0000010000011100_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6613] = 33'b0000110000011100_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6614] = 33'b0000110000011100_0_0_00_000_000_000_0_0_00;
      patterns[6615] = 33'b1000010001110011_0_1_00_111_011_100_0_x_00;
      patterns[6616] = 33'b1000110001110011_1_1_00_111_011_100_0_x_00;
      patterns[6617] = 33'b1000110001110011_0_0_00_000_000_000_0_0_00;
      patterns[6618] = 33'b1001010001110011_0_1_01_111_011_100_0_x_00;
      patterns[6619] = 33'b1001110001110011_1_1_01_111_011_100_0_x_00;
      patterns[6620] = 33'b1001110001110011_0_0_00_000_000_000_0_0_00;
      patterns[6621] = 33'b1010010001110011_0_1_10_111_011_100_0_x_00;
      patterns[6622] = 33'b1010110001110011_1_1_10_111_011_100_0_x_00;
      patterns[6623] = 33'b1010110001110011_0_0_00_000_000_000_0_0_00;
      patterns[6624] = 33'b1011010001110011_0_1_11_111_011_100_0_x_00;
      patterns[6625] = 33'b1011110001110011_1_1_11_111_011_100_0_x_00;
      patterns[6626] = 33'b1011110001110011_0_0_00_000_000_000_0_0_00;
      patterns[6627] = 33'b0101010001110000_0_1_xx_111_xxx_100_0_1_01;
      patterns[6628] = 33'b0101110001110000_1_1_xx_111_xxx_100_0_1_01;
      patterns[6629] = 33'b0101110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6630] = 33'b0100010001110000_0_0_xx_111_100_xxx_1_x_xx;
      patterns[6631] = 33'b0100110001110000_1_0_xx_111_100_xxx_1_x_xx;
      patterns[6632] = 33'b0100110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6633] = 33'b0000010001000010_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6634] = 33'b0000110001000010_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6635] = 33'b0000110001000010_0_0_00_000_000_000_0_0_00;
      patterns[6636] = 33'b1000010001110100_0_1_00_111_100_100_0_x_00;
      patterns[6637] = 33'b1000110001110100_1_1_00_111_100_100_0_x_00;
      patterns[6638] = 33'b1000110001110100_0_0_00_000_000_000_0_0_00;
      patterns[6639] = 33'b1001010001110100_0_1_01_111_100_100_0_x_00;
      patterns[6640] = 33'b1001110001110100_1_1_01_111_100_100_0_x_00;
      patterns[6641] = 33'b1001110001110100_0_0_00_000_000_000_0_0_00;
      patterns[6642] = 33'b1010010001110100_0_1_10_111_100_100_0_x_00;
      patterns[6643] = 33'b1010110001110100_1_1_10_111_100_100_0_x_00;
      patterns[6644] = 33'b1010110001110100_0_0_00_000_000_000_0_0_00;
      patterns[6645] = 33'b1011010001110100_0_1_11_111_100_100_0_x_00;
      patterns[6646] = 33'b1011110001110100_1_1_11_111_100_100_0_x_00;
      patterns[6647] = 33'b1011110001110100_0_0_00_000_000_000_0_0_00;
      patterns[6648] = 33'b0101010001110000_0_1_xx_111_xxx_100_0_1_01;
      patterns[6649] = 33'b0101110001110000_1_1_xx_111_xxx_100_0_1_01;
      patterns[6650] = 33'b0101110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6651] = 33'b0100010001110000_0_0_xx_111_100_xxx_1_x_xx;
      patterns[6652] = 33'b0100110001110000_1_0_xx_111_100_xxx_1_x_xx;
      patterns[6653] = 33'b0100110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6654] = 33'b0000010011101101_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6655] = 33'b0000110011101101_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6656] = 33'b0000110011101101_0_0_00_000_000_000_0_0_00;
      patterns[6657] = 33'b1000010001110101_0_1_00_111_101_100_0_x_00;
      patterns[6658] = 33'b1000110001110101_1_1_00_111_101_100_0_x_00;
      patterns[6659] = 33'b1000110001110101_0_0_00_000_000_000_0_0_00;
      patterns[6660] = 33'b1001010001110101_0_1_01_111_101_100_0_x_00;
      patterns[6661] = 33'b1001110001110101_1_1_01_111_101_100_0_x_00;
      patterns[6662] = 33'b1001110001110101_0_0_00_000_000_000_0_0_00;
      patterns[6663] = 33'b1010010001110101_0_1_10_111_101_100_0_x_00;
      patterns[6664] = 33'b1010110001110101_1_1_10_111_101_100_0_x_00;
      patterns[6665] = 33'b1010110001110101_0_0_00_000_000_000_0_0_00;
      patterns[6666] = 33'b1011010001110101_0_1_11_111_101_100_0_x_00;
      patterns[6667] = 33'b1011110001110101_1_1_11_111_101_100_0_x_00;
      patterns[6668] = 33'b1011110001110101_0_0_00_000_000_000_0_0_00;
      patterns[6669] = 33'b0101010001110000_0_1_xx_111_xxx_100_0_1_01;
      patterns[6670] = 33'b0101110001110000_1_1_xx_111_xxx_100_0_1_01;
      patterns[6671] = 33'b0101110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6672] = 33'b0100010001110000_0_0_xx_111_100_xxx_1_x_xx;
      patterns[6673] = 33'b0100110001110000_1_0_xx_111_100_xxx_1_x_xx;
      patterns[6674] = 33'b0100110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6675] = 33'b0000010000000001_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6676] = 33'b0000110000000001_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6677] = 33'b0000110000000001_0_0_00_000_000_000_0_0_00;
      patterns[6678] = 33'b1000010001110110_0_1_00_111_110_100_0_x_00;
      patterns[6679] = 33'b1000110001110110_1_1_00_111_110_100_0_x_00;
      patterns[6680] = 33'b1000110001110110_0_0_00_000_000_000_0_0_00;
      patterns[6681] = 33'b1001010001110110_0_1_01_111_110_100_0_x_00;
      patterns[6682] = 33'b1001110001110110_1_1_01_111_110_100_0_x_00;
      patterns[6683] = 33'b1001110001110110_0_0_00_000_000_000_0_0_00;
      patterns[6684] = 33'b1010010001110110_0_1_10_111_110_100_0_x_00;
      patterns[6685] = 33'b1010110001110110_1_1_10_111_110_100_0_x_00;
      patterns[6686] = 33'b1010110001110110_0_0_00_000_000_000_0_0_00;
      patterns[6687] = 33'b1011010001110110_0_1_11_111_110_100_0_x_00;
      patterns[6688] = 33'b1011110001110110_1_1_11_111_110_100_0_x_00;
      patterns[6689] = 33'b1011110001110110_0_0_00_000_000_000_0_0_00;
      patterns[6690] = 33'b0101010001110000_0_1_xx_111_xxx_100_0_1_01;
      patterns[6691] = 33'b0101110001110000_1_1_xx_111_xxx_100_0_1_01;
      patterns[6692] = 33'b0101110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6693] = 33'b0100010001110000_0_0_xx_111_100_xxx_1_x_xx;
      patterns[6694] = 33'b0100110001110000_1_0_xx_111_100_xxx_1_x_xx;
      patterns[6695] = 33'b0100110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6696] = 33'b0000010001100111_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6697] = 33'b0000110001100111_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6698] = 33'b0000110001100111_0_0_00_000_000_000_0_0_00;
      patterns[6699] = 33'b1000010001110111_0_1_00_111_111_100_0_x_00;
      patterns[6700] = 33'b1000110001110111_1_1_00_111_111_100_0_x_00;
      patterns[6701] = 33'b1000110001110111_0_0_00_000_000_000_0_0_00;
      patterns[6702] = 33'b1001010001110111_0_1_01_111_111_100_0_x_00;
      patterns[6703] = 33'b1001110001110111_1_1_01_111_111_100_0_x_00;
      patterns[6704] = 33'b1001110001110111_0_0_00_000_000_000_0_0_00;
      patterns[6705] = 33'b1010010001110111_0_1_10_111_111_100_0_x_00;
      patterns[6706] = 33'b1010110001110111_1_1_10_111_111_100_0_x_00;
      patterns[6707] = 33'b1010110001110111_0_0_00_000_000_000_0_0_00;
      patterns[6708] = 33'b1011010001110111_0_1_11_111_111_100_0_x_00;
      patterns[6709] = 33'b1011110001110111_1_1_11_111_111_100_0_x_00;
      patterns[6710] = 33'b1011110001110111_0_0_00_000_000_000_0_0_00;
      patterns[6711] = 33'b0101010001110000_0_1_xx_111_xxx_100_0_1_01;
      patterns[6712] = 33'b0101110001110000_1_1_xx_111_xxx_100_0_1_01;
      patterns[6713] = 33'b0101110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6714] = 33'b0100010001110000_0_0_xx_111_100_xxx_1_x_xx;
      patterns[6715] = 33'b0100110001110000_1_0_xx_111_100_xxx_1_x_xx;
      patterns[6716] = 33'b0100110001110000_0_0_00_000_000_000_0_0_00;
      patterns[6717] = 33'b0000010000001110_0_1_xx_xxx_xxx_100_0_x_10;
      patterns[6718] = 33'b0000110000001110_1_1_xx_xxx_xxx_100_0_x_10;
      patterns[6719] = 33'b0000110000001110_0_0_00_000_000_000_0_0_00;
      patterns[6720] = 33'b1000010100000000_0_1_00_000_000_101_0_x_00;
      patterns[6721] = 33'b1000110100000000_1_1_00_000_000_101_0_x_00;
      patterns[6722] = 33'b1000110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6723] = 33'b1001010100000000_0_1_01_000_000_101_0_x_00;
      patterns[6724] = 33'b1001110100000000_1_1_01_000_000_101_0_x_00;
      patterns[6725] = 33'b1001110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6726] = 33'b1010010100000000_0_1_10_000_000_101_0_x_00;
      patterns[6727] = 33'b1010110100000000_1_1_10_000_000_101_0_x_00;
      patterns[6728] = 33'b1010110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6729] = 33'b1011010100000000_0_1_11_000_000_101_0_x_00;
      patterns[6730] = 33'b1011110100000000_1_1_11_000_000_101_0_x_00;
      patterns[6731] = 33'b1011110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6732] = 33'b0101010100000000_0_1_xx_000_xxx_101_0_1_01;
      patterns[6733] = 33'b0101110100000000_1_1_xx_000_xxx_101_0_1_01;
      patterns[6734] = 33'b0101110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6735] = 33'b0100010100000000_0_0_xx_000_101_xxx_1_x_xx;
      patterns[6736] = 33'b0100110100000000_1_0_xx_000_101_xxx_1_x_xx;
      patterns[6737] = 33'b0100110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6738] = 33'b0000010111100100_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[6739] = 33'b0000110111100100_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[6740] = 33'b0000110111100100_0_0_00_000_000_000_0_0_00;
      patterns[6741] = 33'b1000010100000001_0_1_00_000_001_101_0_x_00;
      patterns[6742] = 33'b1000110100000001_1_1_00_000_001_101_0_x_00;
      patterns[6743] = 33'b1000110100000001_0_0_00_000_000_000_0_0_00;
      patterns[6744] = 33'b1001010100000001_0_1_01_000_001_101_0_x_00;
      patterns[6745] = 33'b1001110100000001_1_1_01_000_001_101_0_x_00;
      patterns[6746] = 33'b1001110100000001_0_0_00_000_000_000_0_0_00;
      patterns[6747] = 33'b1010010100000001_0_1_10_000_001_101_0_x_00;
      patterns[6748] = 33'b1010110100000001_1_1_10_000_001_101_0_x_00;
      patterns[6749] = 33'b1010110100000001_0_0_00_000_000_000_0_0_00;
      patterns[6750] = 33'b1011010100000001_0_1_11_000_001_101_0_x_00;
      patterns[6751] = 33'b1011110100000001_1_1_11_000_001_101_0_x_00;
      patterns[6752] = 33'b1011110100000001_0_0_00_000_000_000_0_0_00;
      patterns[6753] = 33'b0101010100000000_0_1_xx_000_xxx_101_0_1_01;
      patterns[6754] = 33'b0101110100000000_1_1_xx_000_xxx_101_0_1_01;
      patterns[6755] = 33'b0101110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6756] = 33'b0100010100000000_0_0_xx_000_101_xxx_1_x_xx;
      patterns[6757] = 33'b0100110100000000_1_0_xx_000_101_xxx_1_x_xx;
      patterns[6758] = 33'b0100110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6759] = 33'b0000010111101101_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[6760] = 33'b0000110111101101_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[6761] = 33'b0000110111101101_0_0_00_000_000_000_0_0_00;
      patterns[6762] = 33'b1000010100000010_0_1_00_000_010_101_0_x_00;
      patterns[6763] = 33'b1000110100000010_1_1_00_000_010_101_0_x_00;
      patterns[6764] = 33'b1000110100000010_0_0_00_000_000_000_0_0_00;
      patterns[6765] = 33'b1001010100000010_0_1_01_000_010_101_0_x_00;
      patterns[6766] = 33'b1001110100000010_1_1_01_000_010_101_0_x_00;
      patterns[6767] = 33'b1001110100000010_0_0_00_000_000_000_0_0_00;
      patterns[6768] = 33'b1010010100000010_0_1_10_000_010_101_0_x_00;
      patterns[6769] = 33'b1010110100000010_1_1_10_000_010_101_0_x_00;
      patterns[6770] = 33'b1010110100000010_0_0_00_000_000_000_0_0_00;
      patterns[6771] = 33'b1011010100000010_0_1_11_000_010_101_0_x_00;
      patterns[6772] = 33'b1011110100000010_1_1_11_000_010_101_0_x_00;
      patterns[6773] = 33'b1011110100000010_0_0_00_000_000_000_0_0_00;
      patterns[6774] = 33'b0101010100000000_0_1_xx_000_xxx_101_0_1_01;
      patterns[6775] = 33'b0101110100000000_1_1_xx_000_xxx_101_0_1_01;
      patterns[6776] = 33'b0101110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6777] = 33'b0100010100000000_0_0_xx_000_101_xxx_1_x_xx;
      patterns[6778] = 33'b0100110100000000_1_0_xx_000_101_xxx_1_x_xx;
      patterns[6779] = 33'b0100110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6780] = 33'b0000010101010001_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[6781] = 33'b0000110101010001_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[6782] = 33'b0000110101010001_0_0_00_000_000_000_0_0_00;
      patterns[6783] = 33'b1000010100000011_0_1_00_000_011_101_0_x_00;
      patterns[6784] = 33'b1000110100000011_1_1_00_000_011_101_0_x_00;
      patterns[6785] = 33'b1000110100000011_0_0_00_000_000_000_0_0_00;
      patterns[6786] = 33'b1001010100000011_0_1_01_000_011_101_0_x_00;
      patterns[6787] = 33'b1001110100000011_1_1_01_000_011_101_0_x_00;
      patterns[6788] = 33'b1001110100000011_0_0_00_000_000_000_0_0_00;
      patterns[6789] = 33'b1010010100000011_0_1_10_000_011_101_0_x_00;
      patterns[6790] = 33'b1010110100000011_1_1_10_000_011_101_0_x_00;
      patterns[6791] = 33'b1010110100000011_0_0_00_000_000_000_0_0_00;
      patterns[6792] = 33'b1011010100000011_0_1_11_000_011_101_0_x_00;
      patterns[6793] = 33'b1011110100000011_1_1_11_000_011_101_0_x_00;
      patterns[6794] = 33'b1011110100000011_0_0_00_000_000_000_0_0_00;
      patterns[6795] = 33'b0101010100000000_0_1_xx_000_xxx_101_0_1_01;
      patterns[6796] = 33'b0101110100000000_1_1_xx_000_xxx_101_0_1_01;
      patterns[6797] = 33'b0101110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6798] = 33'b0100010100000000_0_0_xx_000_101_xxx_1_x_xx;
      patterns[6799] = 33'b0100110100000000_1_0_xx_000_101_xxx_1_x_xx;
      patterns[6800] = 33'b0100110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6801] = 33'b0000010100011100_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[6802] = 33'b0000110100011100_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[6803] = 33'b0000110100011100_0_0_00_000_000_000_0_0_00;
      patterns[6804] = 33'b1000010100000100_0_1_00_000_100_101_0_x_00;
      patterns[6805] = 33'b1000110100000100_1_1_00_000_100_101_0_x_00;
      patterns[6806] = 33'b1000110100000100_0_0_00_000_000_000_0_0_00;
      patterns[6807] = 33'b1001010100000100_0_1_01_000_100_101_0_x_00;
      patterns[6808] = 33'b1001110100000100_1_1_01_000_100_101_0_x_00;
      patterns[6809] = 33'b1001110100000100_0_0_00_000_000_000_0_0_00;
      patterns[6810] = 33'b1010010100000100_0_1_10_000_100_101_0_x_00;
      patterns[6811] = 33'b1010110100000100_1_1_10_000_100_101_0_x_00;
      patterns[6812] = 33'b1010110100000100_0_0_00_000_000_000_0_0_00;
      patterns[6813] = 33'b1011010100000100_0_1_11_000_100_101_0_x_00;
      patterns[6814] = 33'b1011110100000100_1_1_11_000_100_101_0_x_00;
      patterns[6815] = 33'b1011110100000100_0_0_00_000_000_000_0_0_00;
      patterns[6816] = 33'b0101010100000000_0_1_xx_000_xxx_101_0_1_01;
      patterns[6817] = 33'b0101110100000000_1_1_xx_000_xxx_101_0_1_01;
      patterns[6818] = 33'b0101110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6819] = 33'b0100010100000000_0_0_xx_000_101_xxx_1_x_xx;
      patterns[6820] = 33'b0100110100000000_1_0_xx_000_101_xxx_1_x_xx;
      patterns[6821] = 33'b0100110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6822] = 33'b0000010100011011_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[6823] = 33'b0000110100011011_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[6824] = 33'b0000110100011011_0_0_00_000_000_000_0_0_00;
      patterns[6825] = 33'b1000010100000101_0_1_00_000_101_101_0_x_00;
      patterns[6826] = 33'b1000110100000101_1_1_00_000_101_101_0_x_00;
      patterns[6827] = 33'b1000110100000101_0_0_00_000_000_000_0_0_00;
      patterns[6828] = 33'b1001010100000101_0_1_01_000_101_101_0_x_00;
      patterns[6829] = 33'b1001110100000101_1_1_01_000_101_101_0_x_00;
      patterns[6830] = 33'b1001110100000101_0_0_00_000_000_000_0_0_00;
      patterns[6831] = 33'b1010010100000101_0_1_10_000_101_101_0_x_00;
      patterns[6832] = 33'b1010110100000101_1_1_10_000_101_101_0_x_00;
      patterns[6833] = 33'b1010110100000101_0_0_00_000_000_000_0_0_00;
      patterns[6834] = 33'b1011010100000101_0_1_11_000_101_101_0_x_00;
      patterns[6835] = 33'b1011110100000101_1_1_11_000_101_101_0_x_00;
      patterns[6836] = 33'b1011110100000101_0_0_00_000_000_000_0_0_00;
      patterns[6837] = 33'b0101010100000000_0_1_xx_000_xxx_101_0_1_01;
      patterns[6838] = 33'b0101110100000000_1_1_xx_000_xxx_101_0_1_01;
      patterns[6839] = 33'b0101110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6840] = 33'b0100010100000000_0_0_xx_000_101_xxx_1_x_xx;
      patterns[6841] = 33'b0100110100000000_1_0_xx_000_101_xxx_1_x_xx;
      patterns[6842] = 33'b0100110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6843] = 33'b0000010110110111_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[6844] = 33'b0000110110110111_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[6845] = 33'b0000110110110111_0_0_00_000_000_000_0_0_00;
      patterns[6846] = 33'b1000010100000110_0_1_00_000_110_101_0_x_00;
      patterns[6847] = 33'b1000110100000110_1_1_00_000_110_101_0_x_00;
      patterns[6848] = 33'b1000110100000110_0_0_00_000_000_000_0_0_00;
      patterns[6849] = 33'b1001010100000110_0_1_01_000_110_101_0_x_00;
      patterns[6850] = 33'b1001110100000110_1_1_01_000_110_101_0_x_00;
      patterns[6851] = 33'b1001110100000110_0_0_00_000_000_000_0_0_00;
      patterns[6852] = 33'b1010010100000110_0_1_10_000_110_101_0_x_00;
      patterns[6853] = 33'b1010110100000110_1_1_10_000_110_101_0_x_00;
      patterns[6854] = 33'b1010110100000110_0_0_00_000_000_000_0_0_00;
      patterns[6855] = 33'b1011010100000110_0_1_11_000_110_101_0_x_00;
      patterns[6856] = 33'b1011110100000110_1_1_11_000_110_101_0_x_00;
      patterns[6857] = 33'b1011110100000110_0_0_00_000_000_000_0_0_00;
      patterns[6858] = 33'b0101010100000000_0_1_xx_000_xxx_101_0_1_01;
      patterns[6859] = 33'b0101110100000000_1_1_xx_000_xxx_101_0_1_01;
      patterns[6860] = 33'b0101110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6861] = 33'b0100010100000000_0_0_xx_000_101_xxx_1_x_xx;
      patterns[6862] = 33'b0100110100000000_1_0_xx_000_101_xxx_1_x_xx;
      patterns[6863] = 33'b0100110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6864] = 33'b0000010101011001_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[6865] = 33'b0000110101011001_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[6866] = 33'b0000110101011001_0_0_00_000_000_000_0_0_00;
      patterns[6867] = 33'b1000010100000111_0_1_00_000_111_101_0_x_00;
      patterns[6868] = 33'b1000110100000111_1_1_00_000_111_101_0_x_00;
      patterns[6869] = 33'b1000110100000111_0_0_00_000_000_000_0_0_00;
      patterns[6870] = 33'b1001010100000111_0_1_01_000_111_101_0_x_00;
      patterns[6871] = 33'b1001110100000111_1_1_01_000_111_101_0_x_00;
      patterns[6872] = 33'b1001110100000111_0_0_00_000_000_000_0_0_00;
      patterns[6873] = 33'b1010010100000111_0_1_10_000_111_101_0_x_00;
      patterns[6874] = 33'b1010110100000111_1_1_10_000_111_101_0_x_00;
      patterns[6875] = 33'b1010110100000111_0_0_00_000_000_000_0_0_00;
      patterns[6876] = 33'b1011010100000111_0_1_11_000_111_101_0_x_00;
      patterns[6877] = 33'b1011110100000111_1_1_11_000_111_101_0_x_00;
      patterns[6878] = 33'b1011110100000111_0_0_00_000_000_000_0_0_00;
      patterns[6879] = 33'b0101010100000000_0_1_xx_000_xxx_101_0_1_01;
      patterns[6880] = 33'b0101110100000000_1_1_xx_000_xxx_101_0_1_01;
      patterns[6881] = 33'b0101110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6882] = 33'b0100010100000000_0_0_xx_000_101_xxx_1_x_xx;
      patterns[6883] = 33'b0100110100000000_1_0_xx_000_101_xxx_1_x_xx;
      patterns[6884] = 33'b0100110100000000_0_0_00_000_000_000_0_0_00;
      patterns[6885] = 33'b0000010111101011_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[6886] = 33'b0000110111101011_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[6887] = 33'b0000110111101011_0_0_00_000_000_000_0_0_00;
      patterns[6888] = 33'b1000010100010000_0_1_00_001_000_101_0_x_00;
      patterns[6889] = 33'b1000110100010000_1_1_00_001_000_101_0_x_00;
      patterns[6890] = 33'b1000110100010000_0_0_00_000_000_000_0_0_00;
      patterns[6891] = 33'b1001010100010000_0_1_01_001_000_101_0_x_00;
      patterns[6892] = 33'b1001110100010000_1_1_01_001_000_101_0_x_00;
      patterns[6893] = 33'b1001110100010000_0_0_00_000_000_000_0_0_00;
      patterns[6894] = 33'b1010010100010000_0_1_10_001_000_101_0_x_00;
      patterns[6895] = 33'b1010110100010000_1_1_10_001_000_101_0_x_00;
      patterns[6896] = 33'b1010110100010000_0_0_00_000_000_000_0_0_00;
      patterns[6897] = 33'b1011010100010000_0_1_11_001_000_101_0_x_00;
      patterns[6898] = 33'b1011110100010000_1_1_11_001_000_101_0_x_00;
      patterns[6899] = 33'b1011110100010000_0_0_00_000_000_000_0_0_00;
      patterns[6900] = 33'b0101010100010000_0_1_xx_001_xxx_101_0_1_01;
      patterns[6901] = 33'b0101110100010000_1_1_xx_001_xxx_101_0_1_01;
      patterns[6902] = 33'b0101110100010000_0_0_00_000_000_000_0_0_00;
      patterns[6903] = 33'b0100010100010000_0_0_xx_001_101_xxx_1_x_xx;
      patterns[6904] = 33'b0100110100010000_1_0_xx_001_101_xxx_1_x_xx;
      patterns[6905] = 33'b0100110100010000_0_0_00_000_000_000_0_0_00;
      patterns[6906] = 33'b0000010111010100_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[6907] = 33'b0000110111010100_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[6908] = 33'b0000110111010100_0_0_00_000_000_000_0_0_00;
      patterns[6909] = 33'b1000010100010001_0_1_00_001_001_101_0_x_00;
      patterns[6910] = 33'b1000110100010001_1_1_00_001_001_101_0_x_00;
      patterns[6911] = 33'b1000110100010001_0_0_00_000_000_000_0_0_00;
      patterns[6912] = 33'b1001010100010001_0_1_01_001_001_101_0_x_00;
      patterns[6913] = 33'b1001110100010001_1_1_01_001_001_101_0_x_00;
      patterns[6914] = 33'b1001110100010001_0_0_00_000_000_000_0_0_00;
      patterns[6915] = 33'b1010010100010001_0_1_10_001_001_101_0_x_00;
      patterns[6916] = 33'b1010110100010001_1_1_10_001_001_101_0_x_00;
      patterns[6917] = 33'b1010110100010001_0_0_00_000_000_000_0_0_00;
      patterns[6918] = 33'b1011010100010001_0_1_11_001_001_101_0_x_00;
      patterns[6919] = 33'b1011110100010001_1_1_11_001_001_101_0_x_00;
      patterns[6920] = 33'b1011110100010001_0_0_00_000_000_000_0_0_00;
      patterns[6921] = 33'b0101010100010000_0_1_xx_001_xxx_101_0_1_01;
      patterns[6922] = 33'b0101110100010000_1_1_xx_001_xxx_101_0_1_01;
      patterns[6923] = 33'b0101110100010000_0_0_00_000_000_000_0_0_00;
      patterns[6924] = 33'b0100010100010000_0_0_xx_001_101_xxx_1_x_xx;
      patterns[6925] = 33'b0100110100010000_1_0_xx_001_101_xxx_1_x_xx;
      patterns[6926] = 33'b0100110100010000_0_0_00_000_000_000_0_0_00;
      patterns[6927] = 33'b0000010100001100_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[6928] = 33'b0000110100001100_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[6929] = 33'b0000110100001100_0_0_00_000_000_000_0_0_00;
      patterns[6930] = 33'b1000010100010010_0_1_00_001_010_101_0_x_00;
      patterns[6931] = 33'b1000110100010010_1_1_00_001_010_101_0_x_00;
      patterns[6932] = 33'b1000110100010010_0_0_00_000_000_000_0_0_00;
      patterns[6933] = 33'b1001010100010010_0_1_01_001_010_101_0_x_00;
      patterns[6934] = 33'b1001110100010010_1_1_01_001_010_101_0_x_00;
      patterns[6935] = 33'b1001110100010010_0_0_00_000_000_000_0_0_00;
      patterns[6936] = 33'b1010010100010010_0_1_10_001_010_101_0_x_00;
      patterns[6937] = 33'b1010110100010010_1_1_10_001_010_101_0_x_00;
      patterns[6938] = 33'b1010110100010010_0_0_00_000_000_000_0_0_00;
      patterns[6939] = 33'b1011010100010010_0_1_11_001_010_101_0_x_00;
      patterns[6940] = 33'b1011110100010010_1_1_11_001_010_101_0_x_00;
      patterns[6941] = 33'b1011110100010010_0_0_00_000_000_000_0_0_00;
      patterns[6942] = 33'b0101010100010000_0_1_xx_001_xxx_101_0_1_01;
      patterns[6943] = 33'b0101110100010000_1_1_xx_001_xxx_101_0_1_01;
      patterns[6944] = 33'b0101110100010000_0_0_00_000_000_000_0_0_00;
      patterns[6945] = 33'b0100010100010000_0_0_xx_001_101_xxx_1_x_xx;
      patterns[6946] = 33'b0100110100010000_1_0_xx_001_101_xxx_1_x_xx;
      patterns[6947] = 33'b0100110100010000_0_0_00_000_000_000_0_0_00;
      patterns[6948] = 33'b0000010100011000_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[6949] = 33'b0000110100011000_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[6950] = 33'b0000110100011000_0_0_00_000_000_000_0_0_00;
      patterns[6951] = 33'b1000010100010011_0_1_00_001_011_101_0_x_00;
      patterns[6952] = 33'b1000110100010011_1_1_00_001_011_101_0_x_00;
      patterns[6953] = 33'b1000110100010011_0_0_00_000_000_000_0_0_00;
      patterns[6954] = 33'b1001010100010011_0_1_01_001_011_101_0_x_00;
      patterns[6955] = 33'b1001110100010011_1_1_01_001_011_101_0_x_00;
      patterns[6956] = 33'b1001110100010011_0_0_00_000_000_000_0_0_00;
      patterns[6957] = 33'b1010010100010011_0_1_10_001_011_101_0_x_00;
      patterns[6958] = 33'b1010110100010011_1_1_10_001_011_101_0_x_00;
      patterns[6959] = 33'b1010110100010011_0_0_00_000_000_000_0_0_00;
      patterns[6960] = 33'b1011010100010011_0_1_11_001_011_101_0_x_00;
      patterns[6961] = 33'b1011110100010011_1_1_11_001_011_101_0_x_00;
      patterns[6962] = 33'b1011110100010011_0_0_00_000_000_000_0_0_00;
      patterns[6963] = 33'b0101010100010000_0_1_xx_001_xxx_101_0_1_01;
      patterns[6964] = 33'b0101110100010000_1_1_xx_001_xxx_101_0_1_01;
      patterns[6965] = 33'b0101110100010000_0_0_00_000_000_000_0_0_00;
      patterns[6966] = 33'b0100010100010000_0_0_xx_001_101_xxx_1_x_xx;
      patterns[6967] = 33'b0100110100010000_1_0_xx_001_101_xxx_1_x_xx;
      patterns[6968] = 33'b0100110100010000_0_0_00_000_000_000_0_0_00;
      patterns[6969] = 33'b0000010111001011_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[6970] = 33'b0000110111001011_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[6971] = 33'b0000110111001011_0_0_00_000_000_000_0_0_00;
      patterns[6972] = 33'b1000010100010100_0_1_00_001_100_101_0_x_00;
      patterns[6973] = 33'b1000110100010100_1_1_00_001_100_101_0_x_00;
      patterns[6974] = 33'b1000110100010100_0_0_00_000_000_000_0_0_00;
      patterns[6975] = 33'b1001010100010100_0_1_01_001_100_101_0_x_00;
      patterns[6976] = 33'b1001110100010100_1_1_01_001_100_101_0_x_00;
      patterns[6977] = 33'b1001110100010100_0_0_00_000_000_000_0_0_00;
      patterns[6978] = 33'b1010010100010100_0_1_10_001_100_101_0_x_00;
      patterns[6979] = 33'b1010110100010100_1_1_10_001_100_101_0_x_00;
      patterns[6980] = 33'b1010110100010100_0_0_00_000_000_000_0_0_00;
      patterns[6981] = 33'b1011010100010100_0_1_11_001_100_101_0_x_00;
      patterns[6982] = 33'b1011110100010100_1_1_11_001_100_101_0_x_00;
      patterns[6983] = 33'b1011110100010100_0_0_00_000_000_000_0_0_00;
      patterns[6984] = 33'b0101010100010000_0_1_xx_001_xxx_101_0_1_01;
      patterns[6985] = 33'b0101110100010000_1_1_xx_001_xxx_101_0_1_01;
      patterns[6986] = 33'b0101110100010000_0_0_00_000_000_000_0_0_00;
      patterns[6987] = 33'b0100010100010000_0_0_xx_001_101_xxx_1_x_xx;
      patterns[6988] = 33'b0100110100010000_1_0_xx_001_101_xxx_1_x_xx;
      patterns[6989] = 33'b0100110100010000_0_0_00_000_000_000_0_0_00;
      patterns[6990] = 33'b0000010110111110_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[6991] = 33'b0000110110111110_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[6992] = 33'b0000110110111110_0_0_00_000_000_000_0_0_00;
      patterns[6993] = 33'b1000010100010101_0_1_00_001_101_101_0_x_00;
      patterns[6994] = 33'b1000110100010101_1_1_00_001_101_101_0_x_00;
      patterns[6995] = 33'b1000110100010101_0_0_00_000_000_000_0_0_00;
      patterns[6996] = 33'b1001010100010101_0_1_01_001_101_101_0_x_00;
      patterns[6997] = 33'b1001110100010101_1_1_01_001_101_101_0_x_00;
      patterns[6998] = 33'b1001110100010101_0_0_00_000_000_000_0_0_00;
      patterns[6999] = 33'b1010010100010101_0_1_10_001_101_101_0_x_00;
      patterns[7000] = 33'b1010110100010101_1_1_10_001_101_101_0_x_00;
      patterns[7001] = 33'b1010110100010101_0_0_00_000_000_000_0_0_00;
      patterns[7002] = 33'b1011010100010101_0_1_11_001_101_101_0_x_00;
      patterns[7003] = 33'b1011110100010101_1_1_11_001_101_101_0_x_00;
      patterns[7004] = 33'b1011110100010101_0_0_00_000_000_000_0_0_00;
      patterns[7005] = 33'b0101010100010000_0_1_xx_001_xxx_101_0_1_01;
      patterns[7006] = 33'b0101110100010000_1_1_xx_001_xxx_101_0_1_01;
      patterns[7007] = 33'b0101110100010000_0_0_00_000_000_000_0_0_00;
      patterns[7008] = 33'b0100010100010000_0_0_xx_001_101_xxx_1_x_xx;
      patterns[7009] = 33'b0100110100010000_1_0_xx_001_101_xxx_1_x_xx;
      patterns[7010] = 33'b0100110100010000_0_0_00_000_000_000_0_0_00;
      patterns[7011] = 33'b0000010101001101_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7012] = 33'b0000110101001101_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7013] = 33'b0000110101001101_0_0_00_000_000_000_0_0_00;
      patterns[7014] = 33'b1000010100010110_0_1_00_001_110_101_0_x_00;
      patterns[7015] = 33'b1000110100010110_1_1_00_001_110_101_0_x_00;
      patterns[7016] = 33'b1000110100010110_0_0_00_000_000_000_0_0_00;
      patterns[7017] = 33'b1001010100010110_0_1_01_001_110_101_0_x_00;
      patterns[7018] = 33'b1001110100010110_1_1_01_001_110_101_0_x_00;
      patterns[7019] = 33'b1001110100010110_0_0_00_000_000_000_0_0_00;
      patterns[7020] = 33'b1010010100010110_0_1_10_001_110_101_0_x_00;
      patterns[7021] = 33'b1010110100010110_1_1_10_001_110_101_0_x_00;
      patterns[7022] = 33'b1010110100010110_0_0_00_000_000_000_0_0_00;
      patterns[7023] = 33'b1011010100010110_0_1_11_001_110_101_0_x_00;
      patterns[7024] = 33'b1011110100010110_1_1_11_001_110_101_0_x_00;
      patterns[7025] = 33'b1011110100010110_0_0_00_000_000_000_0_0_00;
      patterns[7026] = 33'b0101010100010000_0_1_xx_001_xxx_101_0_1_01;
      patterns[7027] = 33'b0101110100010000_1_1_xx_001_xxx_101_0_1_01;
      patterns[7028] = 33'b0101110100010000_0_0_00_000_000_000_0_0_00;
      patterns[7029] = 33'b0100010100010000_0_0_xx_001_101_xxx_1_x_xx;
      patterns[7030] = 33'b0100110100010000_1_0_xx_001_101_xxx_1_x_xx;
      patterns[7031] = 33'b0100110100010000_0_0_00_000_000_000_0_0_00;
      patterns[7032] = 33'b0000010100010011_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7033] = 33'b0000110100010011_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7034] = 33'b0000110100010011_0_0_00_000_000_000_0_0_00;
      patterns[7035] = 33'b1000010100010111_0_1_00_001_111_101_0_x_00;
      patterns[7036] = 33'b1000110100010111_1_1_00_001_111_101_0_x_00;
      patterns[7037] = 33'b1000110100010111_0_0_00_000_000_000_0_0_00;
      patterns[7038] = 33'b1001010100010111_0_1_01_001_111_101_0_x_00;
      patterns[7039] = 33'b1001110100010111_1_1_01_001_111_101_0_x_00;
      patterns[7040] = 33'b1001110100010111_0_0_00_000_000_000_0_0_00;
      patterns[7041] = 33'b1010010100010111_0_1_10_001_111_101_0_x_00;
      patterns[7042] = 33'b1010110100010111_1_1_10_001_111_101_0_x_00;
      patterns[7043] = 33'b1010110100010111_0_0_00_000_000_000_0_0_00;
      patterns[7044] = 33'b1011010100010111_0_1_11_001_111_101_0_x_00;
      patterns[7045] = 33'b1011110100010111_1_1_11_001_111_101_0_x_00;
      patterns[7046] = 33'b1011110100010111_0_0_00_000_000_000_0_0_00;
      patterns[7047] = 33'b0101010100010000_0_1_xx_001_xxx_101_0_1_01;
      patterns[7048] = 33'b0101110100010000_1_1_xx_001_xxx_101_0_1_01;
      patterns[7049] = 33'b0101110100010000_0_0_00_000_000_000_0_0_00;
      patterns[7050] = 33'b0100010100010000_0_0_xx_001_101_xxx_1_x_xx;
      patterns[7051] = 33'b0100110100010000_1_0_xx_001_101_xxx_1_x_xx;
      patterns[7052] = 33'b0100110100010000_0_0_00_000_000_000_0_0_00;
      patterns[7053] = 33'b0000010111001110_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7054] = 33'b0000110111001110_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7055] = 33'b0000110111001110_0_0_00_000_000_000_0_0_00;
      patterns[7056] = 33'b1000010100100000_0_1_00_010_000_101_0_x_00;
      patterns[7057] = 33'b1000110100100000_1_1_00_010_000_101_0_x_00;
      patterns[7058] = 33'b1000110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7059] = 33'b1001010100100000_0_1_01_010_000_101_0_x_00;
      patterns[7060] = 33'b1001110100100000_1_1_01_010_000_101_0_x_00;
      patterns[7061] = 33'b1001110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7062] = 33'b1010010100100000_0_1_10_010_000_101_0_x_00;
      patterns[7063] = 33'b1010110100100000_1_1_10_010_000_101_0_x_00;
      patterns[7064] = 33'b1010110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7065] = 33'b1011010100100000_0_1_11_010_000_101_0_x_00;
      patterns[7066] = 33'b1011110100100000_1_1_11_010_000_101_0_x_00;
      patterns[7067] = 33'b1011110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7068] = 33'b0101010100100000_0_1_xx_010_xxx_101_0_1_01;
      patterns[7069] = 33'b0101110100100000_1_1_xx_010_xxx_101_0_1_01;
      patterns[7070] = 33'b0101110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7071] = 33'b0100010100100000_0_0_xx_010_101_xxx_1_x_xx;
      patterns[7072] = 33'b0100110100100000_1_0_xx_010_101_xxx_1_x_xx;
      patterns[7073] = 33'b0100110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7074] = 33'b0000010110110111_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7075] = 33'b0000110110110111_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7076] = 33'b0000110110110111_0_0_00_000_000_000_0_0_00;
      patterns[7077] = 33'b1000010100100001_0_1_00_010_001_101_0_x_00;
      patterns[7078] = 33'b1000110100100001_1_1_00_010_001_101_0_x_00;
      patterns[7079] = 33'b1000110100100001_0_0_00_000_000_000_0_0_00;
      patterns[7080] = 33'b1001010100100001_0_1_01_010_001_101_0_x_00;
      patterns[7081] = 33'b1001110100100001_1_1_01_010_001_101_0_x_00;
      patterns[7082] = 33'b1001110100100001_0_0_00_000_000_000_0_0_00;
      patterns[7083] = 33'b1010010100100001_0_1_10_010_001_101_0_x_00;
      patterns[7084] = 33'b1010110100100001_1_1_10_010_001_101_0_x_00;
      patterns[7085] = 33'b1010110100100001_0_0_00_000_000_000_0_0_00;
      patterns[7086] = 33'b1011010100100001_0_1_11_010_001_101_0_x_00;
      patterns[7087] = 33'b1011110100100001_1_1_11_010_001_101_0_x_00;
      patterns[7088] = 33'b1011110100100001_0_0_00_000_000_000_0_0_00;
      patterns[7089] = 33'b0101010100100000_0_1_xx_010_xxx_101_0_1_01;
      patterns[7090] = 33'b0101110100100000_1_1_xx_010_xxx_101_0_1_01;
      patterns[7091] = 33'b0101110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7092] = 33'b0100010100100000_0_0_xx_010_101_xxx_1_x_xx;
      patterns[7093] = 33'b0100110100100000_1_0_xx_010_101_xxx_1_x_xx;
      patterns[7094] = 33'b0100110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7095] = 33'b0000010110010111_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7096] = 33'b0000110110010111_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7097] = 33'b0000110110010111_0_0_00_000_000_000_0_0_00;
      patterns[7098] = 33'b1000010100100010_0_1_00_010_010_101_0_x_00;
      patterns[7099] = 33'b1000110100100010_1_1_00_010_010_101_0_x_00;
      patterns[7100] = 33'b1000110100100010_0_0_00_000_000_000_0_0_00;
      patterns[7101] = 33'b1001010100100010_0_1_01_010_010_101_0_x_00;
      patterns[7102] = 33'b1001110100100010_1_1_01_010_010_101_0_x_00;
      patterns[7103] = 33'b1001110100100010_0_0_00_000_000_000_0_0_00;
      patterns[7104] = 33'b1010010100100010_0_1_10_010_010_101_0_x_00;
      patterns[7105] = 33'b1010110100100010_1_1_10_010_010_101_0_x_00;
      patterns[7106] = 33'b1010110100100010_0_0_00_000_000_000_0_0_00;
      patterns[7107] = 33'b1011010100100010_0_1_11_010_010_101_0_x_00;
      patterns[7108] = 33'b1011110100100010_1_1_11_010_010_101_0_x_00;
      patterns[7109] = 33'b1011110100100010_0_0_00_000_000_000_0_0_00;
      patterns[7110] = 33'b0101010100100000_0_1_xx_010_xxx_101_0_1_01;
      patterns[7111] = 33'b0101110100100000_1_1_xx_010_xxx_101_0_1_01;
      patterns[7112] = 33'b0101110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7113] = 33'b0100010100100000_0_0_xx_010_101_xxx_1_x_xx;
      patterns[7114] = 33'b0100110100100000_1_0_xx_010_101_xxx_1_x_xx;
      patterns[7115] = 33'b0100110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7116] = 33'b0000010111011000_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7117] = 33'b0000110111011000_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7118] = 33'b0000110111011000_0_0_00_000_000_000_0_0_00;
      patterns[7119] = 33'b1000010100100011_0_1_00_010_011_101_0_x_00;
      patterns[7120] = 33'b1000110100100011_1_1_00_010_011_101_0_x_00;
      patterns[7121] = 33'b1000110100100011_0_0_00_000_000_000_0_0_00;
      patterns[7122] = 33'b1001010100100011_0_1_01_010_011_101_0_x_00;
      patterns[7123] = 33'b1001110100100011_1_1_01_010_011_101_0_x_00;
      patterns[7124] = 33'b1001110100100011_0_0_00_000_000_000_0_0_00;
      patterns[7125] = 33'b1010010100100011_0_1_10_010_011_101_0_x_00;
      patterns[7126] = 33'b1010110100100011_1_1_10_010_011_101_0_x_00;
      patterns[7127] = 33'b1010110100100011_0_0_00_000_000_000_0_0_00;
      patterns[7128] = 33'b1011010100100011_0_1_11_010_011_101_0_x_00;
      patterns[7129] = 33'b1011110100100011_1_1_11_010_011_101_0_x_00;
      patterns[7130] = 33'b1011110100100011_0_0_00_000_000_000_0_0_00;
      patterns[7131] = 33'b0101010100100000_0_1_xx_010_xxx_101_0_1_01;
      patterns[7132] = 33'b0101110100100000_1_1_xx_010_xxx_101_0_1_01;
      patterns[7133] = 33'b0101110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7134] = 33'b0100010100100000_0_0_xx_010_101_xxx_1_x_xx;
      patterns[7135] = 33'b0100110100100000_1_0_xx_010_101_xxx_1_x_xx;
      patterns[7136] = 33'b0100110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7137] = 33'b0000010110000110_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7138] = 33'b0000110110000110_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7139] = 33'b0000110110000110_0_0_00_000_000_000_0_0_00;
      patterns[7140] = 33'b1000010100100100_0_1_00_010_100_101_0_x_00;
      patterns[7141] = 33'b1000110100100100_1_1_00_010_100_101_0_x_00;
      patterns[7142] = 33'b1000110100100100_0_0_00_000_000_000_0_0_00;
      patterns[7143] = 33'b1001010100100100_0_1_01_010_100_101_0_x_00;
      patterns[7144] = 33'b1001110100100100_1_1_01_010_100_101_0_x_00;
      patterns[7145] = 33'b1001110100100100_0_0_00_000_000_000_0_0_00;
      patterns[7146] = 33'b1010010100100100_0_1_10_010_100_101_0_x_00;
      patterns[7147] = 33'b1010110100100100_1_1_10_010_100_101_0_x_00;
      patterns[7148] = 33'b1010110100100100_0_0_00_000_000_000_0_0_00;
      patterns[7149] = 33'b1011010100100100_0_1_11_010_100_101_0_x_00;
      patterns[7150] = 33'b1011110100100100_1_1_11_010_100_101_0_x_00;
      patterns[7151] = 33'b1011110100100100_0_0_00_000_000_000_0_0_00;
      patterns[7152] = 33'b0101010100100000_0_1_xx_010_xxx_101_0_1_01;
      patterns[7153] = 33'b0101110100100000_1_1_xx_010_xxx_101_0_1_01;
      patterns[7154] = 33'b0101110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7155] = 33'b0100010100100000_0_0_xx_010_101_xxx_1_x_xx;
      patterns[7156] = 33'b0100110100100000_1_0_xx_010_101_xxx_1_x_xx;
      patterns[7157] = 33'b0100110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7158] = 33'b0000010100000010_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7159] = 33'b0000110100000010_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7160] = 33'b0000110100000010_0_0_00_000_000_000_0_0_00;
      patterns[7161] = 33'b1000010100100101_0_1_00_010_101_101_0_x_00;
      patterns[7162] = 33'b1000110100100101_1_1_00_010_101_101_0_x_00;
      patterns[7163] = 33'b1000110100100101_0_0_00_000_000_000_0_0_00;
      patterns[7164] = 33'b1001010100100101_0_1_01_010_101_101_0_x_00;
      patterns[7165] = 33'b1001110100100101_1_1_01_010_101_101_0_x_00;
      patterns[7166] = 33'b1001110100100101_0_0_00_000_000_000_0_0_00;
      patterns[7167] = 33'b1010010100100101_0_1_10_010_101_101_0_x_00;
      patterns[7168] = 33'b1010110100100101_1_1_10_010_101_101_0_x_00;
      patterns[7169] = 33'b1010110100100101_0_0_00_000_000_000_0_0_00;
      patterns[7170] = 33'b1011010100100101_0_1_11_010_101_101_0_x_00;
      patterns[7171] = 33'b1011110100100101_1_1_11_010_101_101_0_x_00;
      patterns[7172] = 33'b1011110100100101_0_0_00_000_000_000_0_0_00;
      patterns[7173] = 33'b0101010100100000_0_1_xx_010_xxx_101_0_1_01;
      patterns[7174] = 33'b0101110100100000_1_1_xx_010_xxx_101_0_1_01;
      patterns[7175] = 33'b0101110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7176] = 33'b0100010100100000_0_0_xx_010_101_xxx_1_x_xx;
      patterns[7177] = 33'b0100110100100000_1_0_xx_010_101_xxx_1_x_xx;
      patterns[7178] = 33'b0100110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7179] = 33'b0000010110011111_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7180] = 33'b0000110110011111_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7181] = 33'b0000110110011111_0_0_00_000_000_000_0_0_00;
      patterns[7182] = 33'b1000010100100110_0_1_00_010_110_101_0_x_00;
      patterns[7183] = 33'b1000110100100110_1_1_00_010_110_101_0_x_00;
      patterns[7184] = 33'b1000110100100110_0_0_00_000_000_000_0_0_00;
      patterns[7185] = 33'b1001010100100110_0_1_01_010_110_101_0_x_00;
      patterns[7186] = 33'b1001110100100110_1_1_01_010_110_101_0_x_00;
      patterns[7187] = 33'b1001110100100110_0_0_00_000_000_000_0_0_00;
      patterns[7188] = 33'b1010010100100110_0_1_10_010_110_101_0_x_00;
      patterns[7189] = 33'b1010110100100110_1_1_10_010_110_101_0_x_00;
      patterns[7190] = 33'b1010110100100110_0_0_00_000_000_000_0_0_00;
      patterns[7191] = 33'b1011010100100110_0_1_11_010_110_101_0_x_00;
      patterns[7192] = 33'b1011110100100110_1_1_11_010_110_101_0_x_00;
      patterns[7193] = 33'b1011110100100110_0_0_00_000_000_000_0_0_00;
      patterns[7194] = 33'b0101010100100000_0_1_xx_010_xxx_101_0_1_01;
      patterns[7195] = 33'b0101110100100000_1_1_xx_010_xxx_101_0_1_01;
      patterns[7196] = 33'b0101110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7197] = 33'b0100010100100000_0_0_xx_010_101_xxx_1_x_xx;
      patterns[7198] = 33'b0100110100100000_1_0_xx_010_101_xxx_1_x_xx;
      patterns[7199] = 33'b0100110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7200] = 33'b0000010101011011_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7201] = 33'b0000110101011011_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7202] = 33'b0000110101011011_0_0_00_000_000_000_0_0_00;
      patterns[7203] = 33'b1000010100100111_0_1_00_010_111_101_0_x_00;
      patterns[7204] = 33'b1000110100100111_1_1_00_010_111_101_0_x_00;
      patterns[7205] = 33'b1000110100100111_0_0_00_000_000_000_0_0_00;
      patterns[7206] = 33'b1001010100100111_0_1_01_010_111_101_0_x_00;
      patterns[7207] = 33'b1001110100100111_1_1_01_010_111_101_0_x_00;
      patterns[7208] = 33'b1001110100100111_0_0_00_000_000_000_0_0_00;
      patterns[7209] = 33'b1010010100100111_0_1_10_010_111_101_0_x_00;
      patterns[7210] = 33'b1010110100100111_1_1_10_010_111_101_0_x_00;
      patterns[7211] = 33'b1010110100100111_0_0_00_000_000_000_0_0_00;
      patterns[7212] = 33'b1011010100100111_0_1_11_010_111_101_0_x_00;
      patterns[7213] = 33'b1011110100100111_1_1_11_010_111_101_0_x_00;
      patterns[7214] = 33'b1011110100100111_0_0_00_000_000_000_0_0_00;
      patterns[7215] = 33'b0101010100100000_0_1_xx_010_xxx_101_0_1_01;
      patterns[7216] = 33'b0101110100100000_1_1_xx_010_xxx_101_0_1_01;
      patterns[7217] = 33'b0101110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7218] = 33'b0100010100100000_0_0_xx_010_101_xxx_1_x_xx;
      patterns[7219] = 33'b0100110100100000_1_0_xx_010_101_xxx_1_x_xx;
      patterns[7220] = 33'b0100110100100000_0_0_00_000_000_000_0_0_00;
      patterns[7221] = 33'b0000010110101110_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7222] = 33'b0000110110101110_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7223] = 33'b0000110110101110_0_0_00_000_000_000_0_0_00;
      patterns[7224] = 33'b1000010100110000_0_1_00_011_000_101_0_x_00;
      patterns[7225] = 33'b1000110100110000_1_1_00_011_000_101_0_x_00;
      patterns[7226] = 33'b1000110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7227] = 33'b1001010100110000_0_1_01_011_000_101_0_x_00;
      patterns[7228] = 33'b1001110100110000_1_1_01_011_000_101_0_x_00;
      patterns[7229] = 33'b1001110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7230] = 33'b1010010100110000_0_1_10_011_000_101_0_x_00;
      patterns[7231] = 33'b1010110100110000_1_1_10_011_000_101_0_x_00;
      patterns[7232] = 33'b1010110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7233] = 33'b1011010100110000_0_1_11_011_000_101_0_x_00;
      patterns[7234] = 33'b1011110100110000_1_1_11_011_000_101_0_x_00;
      patterns[7235] = 33'b1011110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7236] = 33'b0101010100110000_0_1_xx_011_xxx_101_0_1_01;
      patterns[7237] = 33'b0101110100110000_1_1_xx_011_xxx_101_0_1_01;
      patterns[7238] = 33'b0101110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7239] = 33'b0100010100110000_0_0_xx_011_101_xxx_1_x_xx;
      patterns[7240] = 33'b0100110100110000_1_0_xx_011_101_xxx_1_x_xx;
      patterns[7241] = 33'b0100110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7242] = 33'b0000010101000100_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7243] = 33'b0000110101000100_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7244] = 33'b0000110101000100_0_0_00_000_000_000_0_0_00;
      patterns[7245] = 33'b1000010100110001_0_1_00_011_001_101_0_x_00;
      patterns[7246] = 33'b1000110100110001_1_1_00_011_001_101_0_x_00;
      patterns[7247] = 33'b1000110100110001_0_0_00_000_000_000_0_0_00;
      patterns[7248] = 33'b1001010100110001_0_1_01_011_001_101_0_x_00;
      patterns[7249] = 33'b1001110100110001_1_1_01_011_001_101_0_x_00;
      patterns[7250] = 33'b1001110100110001_0_0_00_000_000_000_0_0_00;
      patterns[7251] = 33'b1010010100110001_0_1_10_011_001_101_0_x_00;
      patterns[7252] = 33'b1010110100110001_1_1_10_011_001_101_0_x_00;
      patterns[7253] = 33'b1010110100110001_0_0_00_000_000_000_0_0_00;
      patterns[7254] = 33'b1011010100110001_0_1_11_011_001_101_0_x_00;
      patterns[7255] = 33'b1011110100110001_1_1_11_011_001_101_0_x_00;
      patterns[7256] = 33'b1011110100110001_0_0_00_000_000_000_0_0_00;
      patterns[7257] = 33'b0101010100110000_0_1_xx_011_xxx_101_0_1_01;
      patterns[7258] = 33'b0101110100110000_1_1_xx_011_xxx_101_0_1_01;
      patterns[7259] = 33'b0101110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7260] = 33'b0100010100110000_0_0_xx_011_101_xxx_1_x_xx;
      patterns[7261] = 33'b0100110100110000_1_0_xx_011_101_xxx_1_x_xx;
      patterns[7262] = 33'b0100110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7263] = 33'b0000010101011110_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7264] = 33'b0000110101011110_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7265] = 33'b0000110101011110_0_0_00_000_000_000_0_0_00;
      patterns[7266] = 33'b1000010100110010_0_1_00_011_010_101_0_x_00;
      patterns[7267] = 33'b1000110100110010_1_1_00_011_010_101_0_x_00;
      patterns[7268] = 33'b1000110100110010_0_0_00_000_000_000_0_0_00;
      patterns[7269] = 33'b1001010100110010_0_1_01_011_010_101_0_x_00;
      patterns[7270] = 33'b1001110100110010_1_1_01_011_010_101_0_x_00;
      patterns[7271] = 33'b1001110100110010_0_0_00_000_000_000_0_0_00;
      patterns[7272] = 33'b1010010100110010_0_1_10_011_010_101_0_x_00;
      patterns[7273] = 33'b1010110100110010_1_1_10_011_010_101_0_x_00;
      patterns[7274] = 33'b1010110100110010_0_0_00_000_000_000_0_0_00;
      patterns[7275] = 33'b1011010100110010_0_1_11_011_010_101_0_x_00;
      patterns[7276] = 33'b1011110100110010_1_1_11_011_010_101_0_x_00;
      patterns[7277] = 33'b1011110100110010_0_0_00_000_000_000_0_0_00;
      patterns[7278] = 33'b0101010100110000_0_1_xx_011_xxx_101_0_1_01;
      patterns[7279] = 33'b0101110100110000_1_1_xx_011_xxx_101_0_1_01;
      patterns[7280] = 33'b0101110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7281] = 33'b0100010100110000_0_0_xx_011_101_xxx_1_x_xx;
      patterns[7282] = 33'b0100110100110000_1_0_xx_011_101_xxx_1_x_xx;
      patterns[7283] = 33'b0100110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7284] = 33'b0000010110100011_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7285] = 33'b0000110110100011_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7286] = 33'b0000110110100011_0_0_00_000_000_000_0_0_00;
      patterns[7287] = 33'b1000010100110011_0_1_00_011_011_101_0_x_00;
      patterns[7288] = 33'b1000110100110011_1_1_00_011_011_101_0_x_00;
      patterns[7289] = 33'b1000110100110011_0_0_00_000_000_000_0_0_00;
      patterns[7290] = 33'b1001010100110011_0_1_01_011_011_101_0_x_00;
      patterns[7291] = 33'b1001110100110011_1_1_01_011_011_101_0_x_00;
      patterns[7292] = 33'b1001110100110011_0_0_00_000_000_000_0_0_00;
      patterns[7293] = 33'b1010010100110011_0_1_10_011_011_101_0_x_00;
      patterns[7294] = 33'b1010110100110011_1_1_10_011_011_101_0_x_00;
      patterns[7295] = 33'b1010110100110011_0_0_00_000_000_000_0_0_00;
      patterns[7296] = 33'b1011010100110011_0_1_11_011_011_101_0_x_00;
      patterns[7297] = 33'b1011110100110011_1_1_11_011_011_101_0_x_00;
      patterns[7298] = 33'b1011110100110011_0_0_00_000_000_000_0_0_00;
      patterns[7299] = 33'b0101010100110000_0_1_xx_011_xxx_101_0_1_01;
      patterns[7300] = 33'b0101110100110000_1_1_xx_011_xxx_101_0_1_01;
      patterns[7301] = 33'b0101110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7302] = 33'b0100010100110000_0_0_xx_011_101_xxx_1_x_xx;
      patterns[7303] = 33'b0100110100110000_1_0_xx_011_101_xxx_1_x_xx;
      patterns[7304] = 33'b0100110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7305] = 33'b0000010110111000_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7306] = 33'b0000110110111000_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7307] = 33'b0000110110111000_0_0_00_000_000_000_0_0_00;
      patterns[7308] = 33'b1000010100110100_0_1_00_011_100_101_0_x_00;
      patterns[7309] = 33'b1000110100110100_1_1_00_011_100_101_0_x_00;
      patterns[7310] = 33'b1000110100110100_0_0_00_000_000_000_0_0_00;
      patterns[7311] = 33'b1001010100110100_0_1_01_011_100_101_0_x_00;
      patterns[7312] = 33'b1001110100110100_1_1_01_011_100_101_0_x_00;
      patterns[7313] = 33'b1001110100110100_0_0_00_000_000_000_0_0_00;
      patterns[7314] = 33'b1010010100110100_0_1_10_011_100_101_0_x_00;
      patterns[7315] = 33'b1010110100110100_1_1_10_011_100_101_0_x_00;
      patterns[7316] = 33'b1010110100110100_0_0_00_000_000_000_0_0_00;
      patterns[7317] = 33'b1011010100110100_0_1_11_011_100_101_0_x_00;
      patterns[7318] = 33'b1011110100110100_1_1_11_011_100_101_0_x_00;
      patterns[7319] = 33'b1011110100110100_0_0_00_000_000_000_0_0_00;
      patterns[7320] = 33'b0101010100110000_0_1_xx_011_xxx_101_0_1_01;
      patterns[7321] = 33'b0101110100110000_1_1_xx_011_xxx_101_0_1_01;
      patterns[7322] = 33'b0101110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7323] = 33'b0100010100110000_0_0_xx_011_101_xxx_1_x_xx;
      patterns[7324] = 33'b0100110100110000_1_0_xx_011_101_xxx_1_x_xx;
      patterns[7325] = 33'b0100110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7326] = 33'b0000010111101110_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7327] = 33'b0000110111101110_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7328] = 33'b0000110111101110_0_0_00_000_000_000_0_0_00;
      patterns[7329] = 33'b1000010100110101_0_1_00_011_101_101_0_x_00;
      patterns[7330] = 33'b1000110100110101_1_1_00_011_101_101_0_x_00;
      patterns[7331] = 33'b1000110100110101_0_0_00_000_000_000_0_0_00;
      patterns[7332] = 33'b1001010100110101_0_1_01_011_101_101_0_x_00;
      patterns[7333] = 33'b1001110100110101_1_1_01_011_101_101_0_x_00;
      patterns[7334] = 33'b1001110100110101_0_0_00_000_000_000_0_0_00;
      patterns[7335] = 33'b1010010100110101_0_1_10_011_101_101_0_x_00;
      patterns[7336] = 33'b1010110100110101_1_1_10_011_101_101_0_x_00;
      patterns[7337] = 33'b1010110100110101_0_0_00_000_000_000_0_0_00;
      patterns[7338] = 33'b1011010100110101_0_1_11_011_101_101_0_x_00;
      patterns[7339] = 33'b1011110100110101_1_1_11_011_101_101_0_x_00;
      patterns[7340] = 33'b1011110100110101_0_0_00_000_000_000_0_0_00;
      patterns[7341] = 33'b0101010100110000_0_1_xx_011_xxx_101_0_1_01;
      patterns[7342] = 33'b0101110100110000_1_1_xx_011_xxx_101_0_1_01;
      patterns[7343] = 33'b0101110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7344] = 33'b0100010100110000_0_0_xx_011_101_xxx_1_x_xx;
      patterns[7345] = 33'b0100110100110000_1_0_xx_011_101_xxx_1_x_xx;
      patterns[7346] = 33'b0100110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7347] = 33'b0000010110100000_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7348] = 33'b0000110110100000_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7349] = 33'b0000110110100000_0_0_00_000_000_000_0_0_00;
      patterns[7350] = 33'b1000010100110110_0_1_00_011_110_101_0_x_00;
      patterns[7351] = 33'b1000110100110110_1_1_00_011_110_101_0_x_00;
      patterns[7352] = 33'b1000110100110110_0_0_00_000_000_000_0_0_00;
      patterns[7353] = 33'b1001010100110110_0_1_01_011_110_101_0_x_00;
      patterns[7354] = 33'b1001110100110110_1_1_01_011_110_101_0_x_00;
      patterns[7355] = 33'b1001110100110110_0_0_00_000_000_000_0_0_00;
      patterns[7356] = 33'b1010010100110110_0_1_10_011_110_101_0_x_00;
      patterns[7357] = 33'b1010110100110110_1_1_10_011_110_101_0_x_00;
      patterns[7358] = 33'b1010110100110110_0_0_00_000_000_000_0_0_00;
      patterns[7359] = 33'b1011010100110110_0_1_11_011_110_101_0_x_00;
      patterns[7360] = 33'b1011110100110110_1_1_11_011_110_101_0_x_00;
      patterns[7361] = 33'b1011110100110110_0_0_00_000_000_000_0_0_00;
      patterns[7362] = 33'b0101010100110000_0_1_xx_011_xxx_101_0_1_01;
      patterns[7363] = 33'b0101110100110000_1_1_xx_011_xxx_101_0_1_01;
      patterns[7364] = 33'b0101110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7365] = 33'b0100010100110000_0_0_xx_011_101_xxx_1_x_xx;
      patterns[7366] = 33'b0100110100110000_1_0_xx_011_101_xxx_1_x_xx;
      patterns[7367] = 33'b0100110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7368] = 33'b0000010111101100_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7369] = 33'b0000110111101100_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7370] = 33'b0000110111101100_0_0_00_000_000_000_0_0_00;
      patterns[7371] = 33'b1000010100110111_0_1_00_011_111_101_0_x_00;
      patterns[7372] = 33'b1000110100110111_1_1_00_011_111_101_0_x_00;
      patterns[7373] = 33'b1000110100110111_0_0_00_000_000_000_0_0_00;
      patterns[7374] = 33'b1001010100110111_0_1_01_011_111_101_0_x_00;
      patterns[7375] = 33'b1001110100110111_1_1_01_011_111_101_0_x_00;
      patterns[7376] = 33'b1001110100110111_0_0_00_000_000_000_0_0_00;
      patterns[7377] = 33'b1010010100110111_0_1_10_011_111_101_0_x_00;
      patterns[7378] = 33'b1010110100110111_1_1_10_011_111_101_0_x_00;
      patterns[7379] = 33'b1010110100110111_0_0_00_000_000_000_0_0_00;
      patterns[7380] = 33'b1011010100110111_0_1_11_011_111_101_0_x_00;
      patterns[7381] = 33'b1011110100110111_1_1_11_011_111_101_0_x_00;
      patterns[7382] = 33'b1011110100110111_0_0_00_000_000_000_0_0_00;
      patterns[7383] = 33'b0101010100110000_0_1_xx_011_xxx_101_0_1_01;
      patterns[7384] = 33'b0101110100110000_1_1_xx_011_xxx_101_0_1_01;
      patterns[7385] = 33'b0101110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7386] = 33'b0100010100110000_0_0_xx_011_101_xxx_1_x_xx;
      patterns[7387] = 33'b0100110100110000_1_0_xx_011_101_xxx_1_x_xx;
      patterns[7388] = 33'b0100110100110000_0_0_00_000_000_000_0_0_00;
      patterns[7389] = 33'b0000010101100100_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7390] = 33'b0000110101100100_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7391] = 33'b0000110101100100_0_0_00_000_000_000_0_0_00;
      patterns[7392] = 33'b1000010101000000_0_1_00_100_000_101_0_x_00;
      patterns[7393] = 33'b1000110101000000_1_1_00_100_000_101_0_x_00;
      patterns[7394] = 33'b1000110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7395] = 33'b1001010101000000_0_1_01_100_000_101_0_x_00;
      patterns[7396] = 33'b1001110101000000_1_1_01_100_000_101_0_x_00;
      patterns[7397] = 33'b1001110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7398] = 33'b1010010101000000_0_1_10_100_000_101_0_x_00;
      patterns[7399] = 33'b1010110101000000_1_1_10_100_000_101_0_x_00;
      patterns[7400] = 33'b1010110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7401] = 33'b1011010101000000_0_1_11_100_000_101_0_x_00;
      patterns[7402] = 33'b1011110101000000_1_1_11_100_000_101_0_x_00;
      patterns[7403] = 33'b1011110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7404] = 33'b0101010101000000_0_1_xx_100_xxx_101_0_1_01;
      patterns[7405] = 33'b0101110101000000_1_1_xx_100_xxx_101_0_1_01;
      patterns[7406] = 33'b0101110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7407] = 33'b0100010101000000_0_0_xx_100_101_xxx_1_x_xx;
      patterns[7408] = 33'b0100110101000000_1_0_xx_100_101_xxx_1_x_xx;
      patterns[7409] = 33'b0100110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7410] = 33'b0000010101110011_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7411] = 33'b0000110101110011_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7412] = 33'b0000110101110011_0_0_00_000_000_000_0_0_00;
      patterns[7413] = 33'b1000010101000001_0_1_00_100_001_101_0_x_00;
      patterns[7414] = 33'b1000110101000001_1_1_00_100_001_101_0_x_00;
      patterns[7415] = 33'b1000110101000001_0_0_00_000_000_000_0_0_00;
      patterns[7416] = 33'b1001010101000001_0_1_01_100_001_101_0_x_00;
      patterns[7417] = 33'b1001110101000001_1_1_01_100_001_101_0_x_00;
      patterns[7418] = 33'b1001110101000001_0_0_00_000_000_000_0_0_00;
      patterns[7419] = 33'b1010010101000001_0_1_10_100_001_101_0_x_00;
      patterns[7420] = 33'b1010110101000001_1_1_10_100_001_101_0_x_00;
      patterns[7421] = 33'b1010110101000001_0_0_00_000_000_000_0_0_00;
      patterns[7422] = 33'b1011010101000001_0_1_11_100_001_101_0_x_00;
      patterns[7423] = 33'b1011110101000001_1_1_11_100_001_101_0_x_00;
      patterns[7424] = 33'b1011110101000001_0_0_00_000_000_000_0_0_00;
      patterns[7425] = 33'b0101010101000000_0_1_xx_100_xxx_101_0_1_01;
      patterns[7426] = 33'b0101110101000000_1_1_xx_100_xxx_101_0_1_01;
      patterns[7427] = 33'b0101110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7428] = 33'b0100010101000000_0_0_xx_100_101_xxx_1_x_xx;
      patterns[7429] = 33'b0100110101000000_1_0_xx_100_101_xxx_1_x_xx;
      patterns[7430] = 33'b0100110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7431] = 33'b0000010111001110_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7432] = 33'b0000110111001110_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7433] = 33'b0000110111001110_0_0_00_000_000_000_0_0_00;
      patterns[7434] = 33'b1000010101000010_0_1_00_100_010_101_0_x_00;
      patterns[7435] = 33'b1000110101000010_1_1_00_100_010_101_0_x_00;
      patterns[7436] = 33'b1000110101000010_0_0_00_000_000_000_0_0_00;
      patterns[7437] = 33'b1001010101000010_0_1_01_100_010_101_0_x_00;
      patterns[7438] = 33'b1001110101000010_1_1_01_100_010_101_0_x_00;
      patterns[7439] = 33'b1001110101000010_0_0_00_000_000_000_0_0_00;
      patterns[7440] = 33'b1010010101000010_0_1_10_100_010_101_0_x_00;
      patterns[7441] = 33'b1010110101000010_1_1_10_100_010_101_0_x_00;
      patterns[7442] = 33'b1010110101000010_0_0_00_000_000_000_0_0_00;
      patterns[7443] = 33'b1011010101000010_0_1_11_100_010_101_0_x_00;
      patterns[7444] = 33'b1011110101000010_1_1_11_100_010_101_0_x_00;
      patterns[7445] = 33'b1011110101000010_0_0_00_000_000_000_0_0_00;
      patterns[7446] = 33'b0101010101000000_0_1_xx_100_xxx_101_0_1_01;
      patterns[7447] = 33'b0101110101000000_1_1_xx_100_xxx_101_0_1_01;
      patterns[7448] = 33'b0101110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7449] = 33'b0100010101000000_0_0_xx_100_101_xxx_1_x_xx;
      patterns[7450] = 33'b0100110101000000_1_0_xx_100_101_xxx_1_x_xx;
      patterns[7451] = 33'b0100110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7452] = 33'b0000010111110010_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7453] = 33'b0000110111110010_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7454] = 33'b0000110111110010_0_0_00_000_000_000_0_0_00;
      patterns[7455] = 33'b1000010101000011_0_1_00_100_011_101_0_x_00;
      patterns[7456] = 33'b1000110101000011_1_1_00_100_011_101_0_x_00;
      patterns[7457] = 33'b1000110101000011_0_0_00_000_000_000_0_0_00;
      patterns[7458] = 33'b1001010101000011_0_1_01_100_011_101_0_x_00;
      patterns[7459] = 33'b1001110101000011_1_1_01_100_011_101_0_x_00;
      patterns[7460] = 33'b1001110101000011_0_0_00_000_000_000_0_0_00;
      patterns[7461] = 33'b1010010101000011_0_1_10_100_011_101_0_x_00;
      patterns[7462] = 33'b1010110101000011_1_1_10_100_011_101_0_x_00;
      patterns[7463] = 33'b1010110101000011_0_0_00_000_000_000_0_0_00;
      patterns[7464] = 33'b1011010101000011_0_1_11_100_011_101_0_x_00;
      patterns[7465] = 33'b1011110101000011_1_1_11_100_011_101_0_x_00;
      patterns[7466] = 33'b1011110101000011_0_0_00_000_000_000_0_0_00;
      patterns[7467] = 33'b0101010101000000_0_1_xx_100_xxx_101_0_1_01;
      patterns[7468] = 33'b0101110101000000_1_1_xx_100_xxx_101_0_1_01;
      patterns[7469] = 33'b0101110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7470] = 33'b0100010101000000_0_0_xx_100_101_xxx_1_x_xx;
      patterns[7471] = 33'b0100110101000000_1_0_xx_100_101_xxx_1_x_xx;
      patterns[7472] = 33'b0100110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7473] = 33'b0000010101101011_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7474] = 33'b0000110101101011_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7475] = 33'b0000110101101011_0_0_00_000_000_000_0_0_00;
      patterns[7476] = 33'b1000010101000100_0_1_00_100_100_101_0_x_00;
      patterns[7477] = 33'b1000110101000100_1_1_00_100_100_101_0_x_00;
      patterns[7478] = 33'b1000110101000100_0_0_00_000_000_000_0_0_00;
      patterns[7479] = 33'b1001010101000100_0_1_01_100_100_101_0_x_00;
      patterns[7480] = 33'b1001110101000100_1_1_01_100_100_101_0_x_00;
      patterns[7481] = 33'b1001110101000100_0_0_00_000_000_000_0_0_00;
      patterns[7482] = 33'b1010010101000100_0_1_10_100_100_101_0_x_00;
      patterns[7483] = 33'b1010110101000100_1_1_10_100_100_101_0_x_00;
      patterns[7484] = 33'b1010110101000100_0_0_00_000_000_000_0_0_00;
      patterns[7485] = 33'b1011010101000100_0_1_11_100_100_101_0_x_00;
      patterns[7486] = 33'b1011110101000100_1_1_11_100_100_101_0_x_00;
      patterns[7487] = 33'b1011110101000100_0_0_00_000_000_000_0_0_00;
      patterns[7488] = 33'b0101010101000000_0_1_xx_100_xxx_101_0_1_01;
      patterns[7489] = 33'b0101110101000000_1_1_xx_100_xxx_101_0_1_01;
      patterns[7490] = 33'b0101110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7491] = 33'b0100010101000000_0_0_xx_100_101_xxx_1_x_xx;
      patterns[7492] = 33'b0100110101000000_1_0_xx_100_101_xxx_1_x_xx;
      patterns[7493] = 33'b0100110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7494] = 33'b0000010110101010_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7495] = 33'b0000110110101010_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7496] = 33'b0000110110101010_0_0_00_000_000_000_0_0_00;
      patterns[7497] = 33'b1000010101000101_0_1_00_100_101_101_0_x_00;
      patterns[7498] = 33'b1000110101000101_1_1_00_100_101_101_0_x_00;
      patterns[7499] = 33'b1000110101000101_0_0_00_000_000_000_0_0_00;
      patterns[7500] = 33'b1001010101000101_0_1_01_100_101_101_0_x_00;
      patterns[7501] = 33'b1001110101000101_1_1_01_100_101_101_0_x_00;
      patterns[7502] = 33'b1001110101000101_0_0_00_000_000_000_0_0_00;
      patterns[7503] = 33'b1010010101000101_0_1_10_100_101_101_0_x_00;
      patterns[7504] = 33'b1010110101000101_1_1_10_100_101_101_0_x_00;
      patterns[7505] = 33'b1010110101000101_0_0_00_000_000_000_0_0_00;
      patterns[7506] = 33'b1011010101000101_0_1_11_100_101_101_0_x_00;
      patterns[7507] = 33'b1011110101000101_1_1_11_100_101_101_0_x_00;
      patterns[7508] = 33'b1011110101000101_0_0_00_000_000_000_0_0_00;
      patterns[7509] = 33'b0101010101000000_0_1_xx_100_xxx_101_0_1_01;
      patterns[7510] = 33'b0101110101000000_1_1_xx_100_xxx_101_0_1_01;
      patterns[7511] = 33'b0101110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7512] = 33'b0100010101000000_0_0_xx_100_101_xxx_1_x_xx;
      patterns[7513] = 33'b0100110101000000_1_0_xx_100_101_xxx_1_x_xx;
      patterns[7514] = 33'b0100110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7515] = 33'b0000010101101000_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7516] = 33'b0000110101101000_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7517] = 33'b0000110101101000_0_0_00_000_000_000_0_0_00;
      patterns[7518] = 33'b1000010101000110_0_1_00_100_110_101_0_x_00;
      patterns[7519] = 33'b1000110101000110_1_1_00_100_110_101_0_x_00;
      patterns[7520] = 33'b1000110101000110_0_0_00_000_000_000_0_0_00;
      patterns[7521] = 33'b1001010101000110_0_1_01_100_110_101_0_x_00;
      patterns[7522] = 33'b1001110101000110_1_1_01_100_110_101_0_x_00;
      patterns[7523] = 33'b1001110101000110_0_0_00_000_000_000_0_0_00;
      patterns[7524] = 33'b1010010101000110_0_1_10_100_110_101_0_x_00;
      patterns[7525] = 33'b1010110101000110_1_1_10_100_110_101_0_x_00;
      patterns[7526] = 33'b1010110101000110_0_0_00_000_000_000_0_0_00;
      patterns[7527] = 33'b1011010101000110_0_1_11_100_110_101_0_x_00;
      patterns[7528] = 33'b1011110101000110_1_1_11_100_110_101_0_x_00;
      patterns[7529] = 33'b1011110101000110_0_0_00_000_000_000_0_0_00;
      patterns[7530] = 33'b0101010101000000_0_1_xx_100_xxx_101_0_1_01;
      patterns[7531] = 33'b0101110101000000_1_1_xx_100_xxx_101_0_1_01;
      patterns[7532] = 33'b0101110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7533] = 33'b0100010101000000_0_0_xx_100_101_xxx_1_x_xx;
      patterns[7534] = 33'b0100110101000000_1_0_xx_100_101_xxx_1_x_xx;
      patterns[7535] = 33'b0100110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7536] = 33'b0000010110101111_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7537] = 33'b0000110110101111_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7538] = 33'b0000110110101111_0_0_00_000_000_000_0_0_00;
      patterns[7539] = 33'b1000010101000111_0_1_00_100_111_101_0_x_00;
      patterns[7540] = 33'b1000110101000111_1_1_00_100_111_101_0_x_00;
      patterns[7541] = 33'b1000110101000111_0_0_00_000_000_000_0_0_00;
      patterns[7542] = 33'b1001010101000111_0_1_01_100_111_101_0_x_00;
      patterns[7543] = 33'b1001110101000111_1_1_01_100_111_101_0_x_00;
      patterns[7544] = 33'b1001110101000111_0_0_00_000_000_000_0_0_00;
      patterns[7545] = 33'b1010010101000111_0_1_10_100_111_101_0_x_00;
      patterns[7546] = 33'b1010110101000111_1_1_10_100_111_101_0_x_00;
      patterns[7547] = 33'b1010110101000111_0_0_00_000_000_000_0_0_00;
      patterns[7548] = 33'b1011010101000111_0_1_11_100_111_101_0_x_00;
      patterns[7549] = 33'b1011110101000111_1_1_11_100_111_101_0_x_00;
      patterns[7550] = 33'b1011110101000111_0_0_00_000_000_000_0_0_00;
      patterns[7551] = 33'b0101010101000000_0_1_xx_100_xxx_101_0_1_01;
      patterns[7552] = 33'b0101110101000000_1_1_xx_100_xxx_101_0_1_01;
      patterns[7553] = 33'b0101110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7554] = 33'b0100010101000000_0_0_xx_100_101_xxx_1_x_xx;
      patterns[7555] = 33'b0100110101000000_1_0_xx_100_101_xxx_1_x_xx;
      patterns[7556] = 33'b0100110101000000_0_0_00_000_000_000_0_0_00;
      patterns[7557] = 33'b0000010110011110_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7558] = 33'b0000110110011110_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7559] = 33'b0000110110011110_0_0_00_000_000_000_0_0_00;
      patterns[7560] = 33'b1000010101010000_0_1_00_101_000_101_0_x_00;
      patterns[7561] = 33'b1000110101010000_1_1_00_101_000_101_0_x_00;
      patterns[7562] = 33'b1000110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7563] = 33'b1001010101010000_0_1_01_101_000_101_0_x_00;
      patterns[7564] = 33'b1001110101010000_1_1_01_101_000_101_0_x_00;
      patterns[7565] = 33'b1001110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7566] = 33'b1010010101010000_0_1_10_101_000_101_0_x_00;
      patterns[7567] = 33'b1010110101010000_1_1_10_101_000_101_0_x_00;
      patterns[7568] = 33'b1010110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7569] = 33'b1011010101010000_0_1_11_101_000_101_0_x_00;
      patterns[7570] = 33'b1011110101010000_1_1_11_101_000_101_0_x_00;
      patterns[7571] = 33'b1011110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7572] = 33'b0101010101010000_0_1_xx_101_xxx_101_0_1_01;
      patterns[7573] = 33'b0101110101010000_1_1_xx_101_xxx_101_0_1_01;
      patterns[7574] = 33'b0101110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7575] = 33'b0100010101010000_0_0_xx_101_101_xxx_1_x_xx;
      patterns[7576] = 33'b0100110101010000_1_0_xx_101_101_xxx_1_x_xx;
      patterns[7577] = 33'b0100110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7578] = 33'b0000010111111110_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7579] = 33'b0000110111111110_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7580] = 33'b0000110111111110_0_0_00_000_000_000_0_0_00;
      patterns[7581] = 33'b1000010101010001_0_1_00_101_001_101_0_x_00;
      patterns[7582] = 33'b1000110101010001_1_1_00_101_001_101_0_x_00;
      patterns[7583] = 33'b1000110101010001_0_0_00_000_000_000_0_0_00;
      patterns[7584] = 33'b1001010101010001_0_1_01_101_001_101_0_x_00;
      patterns[7585] = 33'b1001110101010001_1_1_01_101_001_101_0_x_00;
      patterns[7586] = 33'b1001110101010001_0_0_00_000_000_000_0_0_00;
      patterns[7587] = 33'b1010010101010001_0_1_10_101_001_101_0_x_00;
      patterns[7588] = 33'b1010110101010001_1_1_10_101_001_101_0_x_00;
      patterns[7589] = 33'b1010110101010001_0_0_00_000_000_000_0_0_00;
      patterns[7590] = 33'b1011010101010001_0_1_11_101_001_101_0_x_00;
      patterns[7591] = 33'b1011110101010001_1_1_11_101_001_101_0_x_00;
      patterns[7592] = 33'b1011110101010001_0_0_00_000_000_000_0_0_00;
      patterns[7593] = 33'b0101010101010000_0_1_xx_101_xxx_101_0_1_01;
      patterns[7594] = 33'b0101110101010000_1_1_xx_101_xxx_101_0_1_01;
      patterns[7595] = 33'b0101110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7596] = 33'b0100010101010000_0_0_xx_101_101_xxx_1_x_xx;
      patterns[7597] = 33'b0100110101010000_1_0_xx_101_101_xxx_1_x_xx;
      patterns[7598] = 33'b0100110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7599] = 33'b0000010111111101_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7600] = 33'b0000110111111101_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7601] = 33'b0000110111111101_0_0_00_000_000_000_0_0_00;
      patterns[7602] = 33'b1000010101010010_0_1_00_101_010_101_0_x_00;
      patterns[7603] = 33'b1000110101010010_1_1_00_101_010_101_0_x_00;
      patterns[7604] = 33'b1000110101010010_0_0_00_000_000_000_0_0_00;
      patterns[7605] = 33'b1001010101010010_0_1_01_101_010_101_0_x_00;
      patterns[7606] = 33'b1001110101010010_1_1_01_101_010_101_0_x_00;
      patterns[7607] = 33'b1001110101010010_0_0_00_000_000_000_0_0_00;
      patterns[7608] = 33'b1010010101010010_0_1_10_101_010_101_0_x_00;
      patterns[7609] = 33'b1010110101010010_1_1_10_101_010_101_0_x_00;
      patterns[7610] = 33'b1010110101010010_0_0_00_000_000_000_0_0_00;
      patterns[7611] = 33'b1011010101010010_0_1_11_101_010_101_0_x_00;
      patterns[7612] = 33'b1011110101010010_1_1_11_101_010_101_0_x_00;
      patterns[7613] = 33'b1011110101010010_0_0_00_000_000_000_0_0_00;
      patterns[7614] = 33'b0101010101010000_0_1_xx_101_xxx_101_0_1_01;
      patterns[7615] = 33'b0101110101010000_1_1_xx_101_xxx_101_0_1_01;
      patterns[7616] = 33'b0101110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7617] = 33'b0100010101010000_0_0_xx_101_101_xxx_1_x_xx;
      patterns[7618] = 33'b0100110101010000_1_0_xx_101_101_xxx_1_x_xx;
      patterns[7619] = 33'b0100110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7620] = 33'b0000010100100101_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7621] = 33'b0000110100100101_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7622] = 33'b0000110100100101_0_0_00_000_000_000_0_0_00;
      patterns[7623] = 33'b1000010101010011_0_1_00_101_011_101_0_x_00;
      patterns[7624] = 33'b1000110101010011_1_1_00_101_011_101_0_x_00;
      patterns[7625] = 33'b1000110101010011_0_0_00_000_000_000_0_0_00;
      patterns[7626] = 33'b1001010101010011_0_1_01_101_011_101_0_x_00;
      patterns[7627] = 33'b1001110101010011_1_1_01_101_011_101_0_x_00;
      patterns[7628] = 33'b1001110101010011_0_0_00_000_000_000_0_0_00;
      patterns[7629] = 33'b1010010101010011_0_1_10_101_011_101_0_x_00;
      patterns[7630] = 33'b1010110101010011_1_1_10_101_011_101_0_x_00;
      patterns[7631] = 33'b1010110101010011_0_0_00_000_000_000_0_0_00;
      patterns[7632] = 33'b1011010101010011_0_1_11_101_011_101_0_x_00;
      patterns[7633] = 33'b1011110101010011_1_1_11_101_011_101_0_x_00;
      patterns[7634] = 33'b1011110101010011_0_0_00_000_000_000_0_0_00;
      patterns[7635] = 33'b0101010101010000_0_1_xx_101_xxx_101_0_1_01;
      patterns[7636] = 33'b0101110101010000_1_1_xx_101_xxx_101_0_1_01;
      patterns[7637] = 33'b0101110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7638] = 33'b0100010101010000_0_0_xx_101_101_xxx_1_x_xx;
      patterns[7639] = 33'b0100110101010000_1_0_xx_101_101_xxx_1_x_xx;
      patterns[7640] = 33'b0100110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7641] = 33'b0000010111000111_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7642] = 33'b0000110111000111_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7643] = 33'b0000110111000111_0_0_00_000_000_000_0_0_00;
      patterns[7644] = 33'b1000010101010100_0_1_00_101_100_101_0_x_00;
      patterns[7645] = 33'b1000110101010100_1_1_00_101_100_101_0_x_00;
      patterns[7646] = 33'b1000110101010100_0_0_00_000_000_000_0_0_00;
      patterns[7647] = 33'b1001010101010100_0_1_01_101_100_101_0_x_00;
      patterns[7648] = 33'b1001110101010100_1_1_01_101_100_101_0_x_00;
      patterns[7649] = 33'b1001110101010100_0_0_00_000_000_000_0_0_00;
      patterns[7650] = 33'b1010010101010100_0_1_10_101_100_101_0_x_00;
      patterns[7651] = 33'b1010110101010100_1_1_10_101_100_101_0_x_00;
      patterns[7652] = 33'b1010110101010100_0_0_00_000_000_000_0_0_00;
      patterns[7653] = 33'b1011010101010100_0_1_11_101_100_101_0_x_00;
      patterns[7654] = 33'b1011110101010100_1_1_11_101_100_101_0_x_00;
      patterns[7655] = 33'b1011110101010100_0_0_00_000_000_000_0_0_00;
      patterns[7656] = 33'b0101010101010000_0_1_xx_101_xxx_101_0_1_01;
      patterns[7657] = 33'b0101110101010000_1_1_xx_101_xxx_101_0_1_01;
      patterns[7658] = 33'b0101110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7659] = 33'b0100010101010000_0_0_xx_101_101_xxx_1_x_xx;
      patterns[7660] = 33'b0100110101010000_1_0_xx_101_101_xxx_1_x_xx;
      patterns[7661] = 33'b0100110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7662] = 33'b0000010110100000_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7663] = 33'b0000110110100000_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7664] = 33'b0000110110100000_0_0_00_000_000_000_0_0_00;
      patterns[7665] = 33'b1000010101010101_0_1_00_101_101_101_0_x_00;
      patterns[7666] = 33'b1000110101010101_1_1_00_101_101_101_0_x_00;
      patterns[7667] = 33'b1000110101010101_0_0_00_000_000_000_0_0_00;
      patterns[7668] = 33'b1001010101010101_0_1_01_101_101_101_0_x_00;
      patterns[7669] = 33'b1001110101010101_1_1_01_101_101_101_0_x_00;
      patterns[7670] = 33'b1001110101010101_0_0_00_000_000_000_0_0_00;
      patterns[7671] = 33'b1010010101010101_0_1_10_101_101_101_0_x_00;
      patterns[7672] = 33'b1010110101010101_1_1_10_101_101_101_0_x_00;
      patterns[7673] = 33'b1010110101010101_0_0_00_000_000_000_0_0_00;
      patterns[7674] = 33'b1011010101010101_0_1_11_101_101_101_0_x_00;
      patterns[7675] = 33'b1011110101010101_1_1_11_101_101_101_0_x_00;
      patterns[7676] = 33'b1011110101010101_0_0_00_000_000_000_0_0_00;
      patterns[7677] = 33'b0101010101010000_0_1_xx_101_xxx_101_0_1_01;
      patterns[7678] = 33'b0101110101010000_1_1_xx_101_xxx_101_0_1_01;
      patterns[7679] = 33'b0101110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7680] = 33'b0100010101010000_0_0_xx_101_101_xxx_1_x_xx;
      patterns[7681] = 33'b0100110101010000_1_0_xx_101_101_xxx_1_x_xx;
      patterns[7682] = 33'b0100110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7683] = 33'b0000010110011011_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7684] = 33'b0000110110011011_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7685] = 33'b0000110110011011_0_0_00_000_000_000_0_0_00;
      patterns[7686] = 33'b1000010101010110_0_1_00_101_110_101_0_x_00;
      patterns[7687] = 33'b1000110101010110_1_1_00_101_110_101_0_x_00;
      patterns[7688] = 33'b1000110101010110_0_0_00_000_000_000_0_0_00;
      patterns[7689] = 33'b1001010101010110_0_1_01_101_110_101_0_x_00;
      patterns[7690] = 33'b1001110101010110_1_1_01_101_110_101_0_x_00;
      patterns[7691] = 33'b1001110101010110_0_0_00_000_000_000_0_0_00;
      patterns[7692] = 33'b1010010101010110_0_1_10_101_110_101_0_x_00;
      patterns[7693] = 33'b1010110101010110_1_1_10_101_110_101_0_x_00;
      patterns[7694] = 33'b1010110101010110_0_0_00_000_000_000_0_0_00;
      patterns[7695] = 33'b1011010101010110_0_1_11_101_110_101_0_x_00;
      patterns[7696] = 33'b1011110101010110_1_1_11_101_110_101_0_x_00;
      patterns[7697] = 33'b1011110101010110_0_0_00_000_000_000_0_0_00;
      patterns[7698] = 33'b0101010101010000_0_1_xx_101_xxx_101_0_1_01;
      patterns[7699] = 33'b0101110101010000_1_1_xx_101_xxx_101_0_1_01;
      patterns[7700] = 33'b0101110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7701] = 33'b0100010101010000_0_0_xx_101_101_xxx_1_x_xx;
      patterns[7702] = 33'b0100110101010000_1_0_xx_101_101_xxx_1_x_xx;
      patterns[7703] = 33'b0100110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7704] = 33'b0000010111001010_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7705] = 33'b0000110111001010_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7706] = 33'b0000110111001010_0_0_00_000_000_000_0_0_00;
      patterns[7707] = 33'b1000010101010111_0_1_00_101_111_101_0_x_00;
      patterns[7708] = 33'b1000110101010111_1_1_00_101_111_101_0_x_00;
      patterns[7709] = 33'b1000110101010111_0_0_00_000_000_000_0_0_00;
      patterns[7710] = 33'b1001010101010111_0_1_01_101_111_101_0_x_00;
      patterns[7711] = 33'b1001110101010111_1_1_01_101_111_101_0_x_00;
      patterns[7712] = 33'b1001110101010111_0_0_00_000_000_000_0_0_00;
      patterns[7713] = 33'b1010010101010111_0_1_10_101_111_101_0_x_00;
      patterns[7714] = 33'b1010110101010111_1_1_10_101_111_101_0_x_00;
      patterns[7715] = 33'b1010110101010111_0_0_00_000_000_000_0_0_00;
      patterns[7716] = 33'b1011010101010111_0_1_11_101_111_101_0_x_00;
      patterns[7717] = 33'b1011110101010111_1_1_11_101_111_101_0_x_00;
      patterns[7718] = 33'b1011110101010111_0_0_00_000_000_000_0_0_00;
      patterns[7719] = 33'b0101010101010000_0_1_xx_101_xxx_101_0_1_01;
      patterns[7720] = 33'b0101110101010000_1_1_xx_101_xxx_101_0_1_01;
      patterns[7721] = 33'b0101110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7722] = 33'b0100010101010000_0_0_xx_101_101_xxx_1_x_xx;
      patterns[7723] = 33'b0100110101010000_1_0_xx_101_101_xxx_1_x_xx;
      patterns[7724] = 33'b0100110101010000_0_0_00_000_000_000_0_0_00;
      patterns[7725] = 33'b0000010111011000_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7726] = 33'b0000110111011000_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7727] = 33'b0000110111011000_0_0_00_000_000_000_0_0_00;
      patterns[7728] = 33'b1000010101100000_0_1_00_110_000_101_0_x_00;
      patterns[7729] = 33'b1000110101100000_1_1_00_110_000_101_0_x_00;
      patterns[7730] = 33'b1000110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7731] = 33'b1001010101100000_0_1_01_110_000_101_0_x_00;
      patterns[7732] = 33'b1001110101100000_1_1_01_110_000_101_0_x_00;
      patterns[7733] = 33'b1001110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7734] = 33'b1010010101100000_0_1_10_110_000_101_0_x_00;
      patterns[7735] = 33'b1010110101100000_1_1_10_110_000_101_0_x_00;
      patterns[7736] = 33'b1010110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7737] = 33'b1011010101100000_0_1_11_110_000_101_0_x_00;
      patterns[7738] = 33'b1011110101100000_1_1_11_110_000_101_0_x_00;
      patterns[7739] = 33'b1011110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7740] = 33'b0101010101100000_0_1_xx_110_xxx_101_0_1_01;
      patterns[7741] = 33'b0101110101100000_1_1_xx_110_xxx_101_0_1_01;
      patterns[7742] = 33'b0101110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7743] = 33'b0100010101100000_0_0_xx_110_101_xxx_1_x_xx;
      patterns[7744] = 33'b0100110101100000_1_0_xx_110_101_xxx_1_x_xx;
      patterns[7745] = 33'b0100110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7746] = 33'b0000010110110010_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7747] = 33'b0000110110110010_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7748] = 33'b0000110110110010_0_0_00_000_000_000_0_0_00;
      patterns[7749] = 33'b1000010101100001_0_1_00_110_001_101_0_x_00;
      patterns[7750] = 33'b1000110101100001_1_1_00_110_001_101_0_x_00;
      patterns[7751] = 33'b1000110101100001_0_0_00_000_000_000_0_0_00;
      patterns[7752] = 33'b1001010101100001_0_1_01_110_001_101_0_x_00;
      patterns[7753] = 33'b1001110101100001_1_1_01_110_001_101_0_x_00;
      patterns[7754] = 33'b1001110101100001_0_0_00_000_000_000_0_0_00;
      patterns[7755] = 33'b1010010101100001_0_1_10_110_001_101_0_x_00;
      patterns[7756] = 33'b1010110101100001_1_1_10_110_001_101_0_x_00;
      patterns[7757] = 33'b1010110101100001_0_0_00_000_000_000_0_0_00;
      patterns[7758] = 33'b1011010101100001_0_1_11_110_001_101_0_x_00;
      patterns[7759] = 33'b1011110101100001_1_1_11_110_001_101_0_x_00;
      patterns[7760] = 33'b1011110101100001_0_0_00_000_000_000_0_0_00;
      patterns[7761] = 33'b0101010101100000_0_1_xx_110_xxx_101_0_1_01;
      patterns[7762] = 33'b0101110101100000_1_1_xx_110_xxx_101_0_1_01;
      patterns[7763] = 33'b0101110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7764] = 33'b0100010101100000_0_0_xx_110_101_xxx_1_x_xx;
      patterns[7765] = 33'b0100110101100000_1_0_xx_110_101_xxx_1_x_xx;
      patterns[7766] = 33'b0100110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7767] = 33'b0000010100011011_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7768] = 33'b0000110100011011_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7769] = 33'b0000110100011011_0_0_00_000_000_000_0_0_00;
      patterns[7770] = 33'b1000010101100010_0_1_00_110_010_101_0_x_00;
      patterns[7771] = 33'b1000110101100010_1_1_00_110_010_101_0_x_00;
      patterns[7772] = 33'b1000110101100010_0_0_00_000_000_000_0_0_00;
      patterns[7773] = 33'b1001010101100010_0_1_01_110_010_101_0_x_00;
      patterns[7774] = 33'b1001110101100010_1_1_01_110_010_101_0_x_00;
      patterns[7775] = 33'b1001110101100010_0_0_00_000_000_000_0_0_00;
      patterns[7776] = 33'b1010010101100010_0_1_10_110_010_101_0_x_00;
      patterns[7777] = 33'b1010110101100010_1_1_10_110_010_101_0_x_00;
      patterns[7778] = 33'b1010110101100010_0_0_00_000_000_000_0_0_00;
      patterns[7779] = 33'b1011010101100010_0_1_11_110_010_101_0_x_00;
      patterns[7780] = 33'b1011110101100010_1_1_11_110_010_101_0_x_00;
      patterns[7781] = 33'b1011110101100010_0_0_00_000_000_000_0_0_00;
      patterns[7782] = 33'b0101010101100000_0_1_xx_110_xxx_101_0_1_01;
      patterns[7783] = 33'b0101110101100000_1_1_xx_110_xxx_101_0_1_01;
      patterns[7784] = 33'b0101110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7785] = 33'b0100010101100000_0_0_xx_110_101_xxx_1_x_xx;
      patterns[7786] = 33'b0100110101100000_1_0_xx_110_101_xxx_1_x_xx;
      patterns[7787] = 33'b0100110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7788] = 33'b0000010100010000_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7789] = 33'b0000110100010000_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7790] = 33'b0000110100010000_0_0_00_000_000_000_0_0_00;
      patterns[7791] = 33'b1000010101100011_0_1_00_110_011_101_0_x_00;
      patterns[7792] = 33'b1000110101100011_1_1_00_110_011_101_0_x_00;
      patterns[7793] = 33'b1000110101100011_0_0_00_000_000_000_0_0_00;
      patterns[7794] = 33'b1001010101100011_0_1_01_110_011_101_0_x_00;
      patterns[7795] = 33'b1001110101100011_1_1_01_110_011_101_0_x_00;
      patterns[7796] = 33'b1001110101100011_0_0_00_000_000_000_0_0_00;
      patterns[7797] = 33'b1010010101100011_0_1_10_110_011_101_0_x_00;
      patterns[7798] = 33'b1010110101100011_1_1_10_110_011_101_0_x_00;
      patterns[7799] = 33'b1010110101100011_0_0_00_000_000_000_0_0_00;
      patterns[7800] = 33'b1011010101100011_0_1_11_110_011_101_0_x_00;
      patterns[7801] = 33'b1011110101100011_1_1_11_110_011_101_0_x_00;
      patterns[7802] = 33'b1011110101100011_0_0_00_000_000_000_0_0_00;
      patterns[7803] = 33'b0101010101100000_0_1_xx_110_xxx_101_0_1_01;
      patterns[7804] = 33'b0101110101100000_1_1_xx_110_xxx_101_0_1_01;
      patterns[7805] = 33'b0101110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7806] = 33'b0100010101100000_0_0_xx_110_101_xxx_1_x_xx;
      patterns[7807] = 33'b0100110101100000_1_0_xx_110_101_xxx_1_x_xx;
      patterns[7808] = 33'b0100110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7809] = 33'b0000010100110111_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7810] = 33'b0000110100110111_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7811] = 33'b0000110100110111_0_0_00_000_000_000_0_0_00;
      patterns[7812] = 33'b1000010101100100_0_1_00_110_100_101_0_x_00;
      patterns[7813] = 33'b1000110101100100_1_1_00_110_100_101_0_x_00;
      patterns[7814] = 33'b1000110101100100_0_0_00_000_000_000_0_0_00;
      patterns[7815] = 33'b1001010101100100_0_1_01_110_100_101_0_x_00;
      patterns[7816] = 33'b1001110101100100_1_1_01_110_100_101_0_x_00;
      patterns[7817] = 33'b1001110101100100_0_0_00_000_000_000_0_0_00;
      patterns[7818] = 33'b1010010101100100_0_1_10_110_100_101_0_x_00;
      patterns[7819] = 33'b1010110101100100_1_1_10_110_100_101_0_x_00;
      patterns[7820] = 33'b1010110101100100_0_0_00_000_000_000_0_0_00;
      patterns[7821] = 33'b1011010101100100_0_1_11_110_100_101_0_x_00;
      patterns[7822] = 33'b1011110101100100_1_1_11_110_100_101_0_x_00;
      patterns[7823] = 33'b1011110101100100_0_0_00_000_000_000_0_0_00;
      patterns[7824] = 33'b0101010101100000_0_1_xx_110_xxx_101_0_1_01;
      patterns[7825] = 33'b0101110101100000_1_1_xx_110_xxx_101_0_1_01;
      patterns[7826] = 33'b0101110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7827] = 33'b0100010101100000_0_0_xx_110_101_xxx_1_x_xx;
      patterns[7828] = 33'b0100110101100000_1_0_xx_110_101_xxx_1_x_xx;
      patterns[7829] = 33'b0100110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7830] = 33'b0000010110001101_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7831] = 33'b0000110110001101_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7832] = 33'b0000110110001101_0_0_00_000_000_000_0_0_00;
      patterns[7833] = 33'b1000010101100101_0_1_00_110_101_101_0_x_00;
      patterns[7834] = 33'b1000110101100101_1_1_00_110_101_101_0_x_00;
      patterns[7835] = 33'b1000110101100101_0_0_00_000_000_000_0_0_00;
      patterns[7836] = 33'b1001010101100101_0_1_01_110_101_101_0_x_00;
      patterns[7837] = 33'b1001110101100101_1_1_01_110_101_101_0_x_00;
      patterns[7838] = 33'b1001110101100101_0_0_00_000_000_000_0_0_00;
      patterns[7839] = 33'b1010010101100101_0_1_10_110_101_101_0_x_00;
      patterns[7840] = 33'b1010110101100101_1_1_10_110_101_101_0_x_00;
      patterns[7841] = 33'b1010110101100101_0_0_00_000_000_000_0_0_00;
      patterns[7842] = 33'b1011010101100101_0_1_11_110_101_101_0_x_00;
      patterns[7843] = 33'b1011110101100101_1_1_11_110_101_101_0_x_00;
      patterns[7844] = 33'b1011110101100101_0_0_00_000_000_000_0_0_00;
      patterns[7845] = 33'b0101010101100000_0_1_xx_110_xxx_101_0_1_01;
      patterns[7846] = 33'b0101110101100000_1_1_xx_110_xxx_101_0_1_01;
      patterns[7847] = 33'b0101110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7848] = 33'b0100010101100000_0_0_xx_110_101_xxx_1_x_xx;
      patterns[7849] = 33'b0100110101100000_1_0_xx_110_101_xxx_1_x_xx;
      patterns[7850] = 33'b0100110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7851] = 33'b0000010111010110_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7852] = 33'b0000110111010110_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7853] = 33'b0000110111010110_0_0_00_000_000_000_0_0_00;
      patterns[7854] = 33'b1000010101100110_0_1_00_110_110_101_0_x_00;
      patterns[7855] = 33'b1000110101100110_1_1_00_110_110_101_0_x_00;
      patterns[7856] = 33'b1000110101100110_0_0_00_000_000_000_0_0_00;
      patterns[7857] = 33'b1001010101100110_0_1_01_110_110_101_0_x_00;
      patterns[7858] = 33'b1001110101100110_1_1_01_110_110_101_0_x_00;
      patterns[7859] = 33'b1001110101100110_0_0_00_000_000_000_0_0_00;
      patterns[7860] = 33'b1010010101100110_0_1_10_110_110_101_0_x_00;
      patterns[7861] = 33'b1010110101100110_1_1_10_110_110_101_0_x_00;
      patterns[7862] = 33'b1010110101100110_0_0_00_000_000_000_0_0_00;
      patterns[7863] = 33'b1011010101100110_0_1_11_110_110_101_0_x_00;
      patterns[7864] = 33'b1011110101100110_1_1_11_110_110_101_0_x_00;
      patterns[7865] = 33'b1011110101100110_0_0_00_000_000_000_0_0_00;
      patterns[7866] = 33'b0101010101100000_0_1_xx_110_xxx_101_0_1_01;
      patterns[7867] = 33'b0101110101100000_1_1_xx_110_xxx_101_0_1_01;
      patterns[7868] = 33'b0101110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7869] = 33'b0100010101100000_0_0_xx_110_101_xxx_1_x_xx;
      patterns[7870] = 33'b0100110101100000_1_0_xx_110_101_xxx_1_x_xx;
      patterns[7871] = 33'b0100110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7872] = 33'b0000010100011111_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7873] = 33'b0000110100011111_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7874] = 33'b0000110100011111_0_0_00_000_000_000_0_0_00;
      patterns[7875] = 33'b1000010101100111_0_1_00_110_111_101_0_x_00;
      patterns[7876] = 33'b1000110101100111_1_1_00_110_111_101_0_x_00;
      patterns[7877] = 33'b1000110101100111_0_0_00_000_000_000_0_0_00;
      patterns[7878] = 33'b1001010101100111_0_1_01_110_111_101_0_x_00;
      patterns[7879] = 33'b1001110101100111_1_1_01_110_111_101_0_x_00;
      patterns[7880] = 33'b1001110101100111_0_0_00_000_000_000_0_0_00;
      patterns[7881] = 33'b1010010101100111_0_1_10_110_111_101_0_x_00;
      patterns[7882] = 33'b1010110101100111_1_1_10_110_111_101_0_x_00;
      patterns[7883] = 33'b1010110101100111_0_0_00_000_000_000_0_0_00;
      patterns[7884] = 33'b1011010101100111_0_1_11_110_111_101_0_x_00;
      patterns[7885] = 33'b1011110101100111_1_1_11_110_111_101_0_x_00;
      patterns[7886] = 33'b1011110101100111_0_0_00_000_000_000_0_0_00;
      patterns[7887] = 33'b0101010101100000_0_1_xx_110_xxx_101_0_1_01;
      patterns[7888] = 33'b0101110101100000_1_1_xx_110_xxx_101_0_1_01;
      patterns[7889] = 33'b0101110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7890] = 33'b0100010101100000_0_0_xx_110_101_xxx_1_x_xx;
      patterns[7891] = 33'b0100110101100000_1_0_xx_110_101_xxx_1_x_xx;
      patterns[7892] = 33'b0100110101100000_0_0_00_000_000_000_0_0_00;
      patterns[7893] = 33'b0000010100001101_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7894] = 33'b0000110100001101_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7895] = 33'b0000110100001101_0_0_00_000_000_000_0_0_00;
      patterns[7896] = 33'b1000010101110000_0_1_00_111_000_101_0_x_00;
      patterns[7897] = 33'b1000110101110000_1_1_00_111_000_101_0_x_00;
      patterns[7898] = 33'b1000110101110000_0_0_00_000_000_000_0_0_00;
      patterns[7899] = 33'b1001010101110000_0_1_01_111_000_101_0_x_00;
      patterns[7900] = 33'b1001110101110000_1_1_01_111_000_101_0_x_00;
      patterns[7901] = 33'b1001110101110000_0_0_00_000_000_000_0_0_00;
      patterns[7902] = 33'b1010010101110000_0_1_10_111_000_101_0_x_00;
      patterns[7903] = 33'b1010110101110000_1_1_10_111_000_101_0_x_00;
      patterns[7904] = 33'b1010110101110000_0_0_00_000_000_000_0_0_00;
      patterns[7905] = 33'b1011010101110000_0_1_11_111_000_101_0_x_00;
      patterns[7906] = 33'b1011110101110000_1_1_11_111_000_101_0_x_00;
      patterns[7907] = 33'b1011110101110000_0_0_00_000_000_000_0_0_00;
      patterns[7908] = 33'b0101010101110000_0_1_xx_111_xxx_101_0_1_01;
      patterns[7909] = 33'b0101110101110000_1_1_xx_111_xxx_101_0_1_01;
      patterns[7910] = 33'b0101110101110000_0_0_00_000_000_000_0_0_00;
      patterns[7911] = 33'b0100010101110000_0_0_xx_111_101_xxx_1_x_xx;
      patterns[7912] = 33'b0100110101110000_1_0_xx_111_101_xxx_1_x_xx;
      patterns[7913] = 33'b0100110101110000_0_0_00_000_000_000_0_0_00;
      patterns[7914] = 33'b0000010110110001_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7915] = 33'b0000110110110001_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7916] = 33'b0000110110110001_0_0_00_000_000_000_0_0_00;
      patterns[7917] = 33'b1000010101110001_0_1_00_111_001_101_0_x_00;
      patterns[7918] = 33'b1000110101110001_1_1_00_111_001_101_0_x_00;
      patterns[7919] = 33'b1000110101110001_0_0_00_000_000_000_0_0_00;
      patterns[7920] = 33'b1001010101110001_0_1_01_111_001_101_0_x_00;
      patterns[7921] = 33'b1001110101110001_1_1_01_111_001_101_0_x_00;
      patterns[7922] = 33'b1001110101110001_0_0_00_000_000_000_0_0_00;
      patterns[7923] = 33'b1010010101110001_0_1_10_111_001_101_0_x_00;
      patterns[7924] = 33'b1010110101110001_1_1_10_111_001_101_0_x_00;
      patterns[7925] = 33'b1010110101110001_0_0_00_000_000_000_0_0_00;
      patterns[7926] = 33'b1011010101110001_0_1_11_111_001_101_0_x_00;
      patterns[7927] = 33'b1011110101110001_1_1_11_111_001_101_0_x_00;
      patterns[7928] = 33'b1011110101110001_0_0_00_000_000_000_0_0_00;
      patterns[7929] = 33'b0101010101110000_0_1_xx_111_xxx_101_0_1_01;
      patterns[7930] = 33'b0101110101110000_1_1_xx_111_xxx_101_0_1_01;
      patterns[7931] = 33'b0101110101110000_0_0_00_000_000_000_0_0_00;
      patterns[7932] = 33'b0100010101110000_0_0_xx_111_101_xxx_1_x_xx;
      patterns[7933] = 33'b0100110101110000_1_0_xx_111_101_xxx_1_x_xx;
      patterns[7934] = 33'b0100110101110000_0_0_00_000_000_000_0_0_00;
      patterns[7935] = 33'b0000010111111110_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7936] = 33'b0000110111111110_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7937] = 33'b0000110111111110_0_0_00_000_000_000_0_0_00;
      patterns[7938] = 33'b1000010101110010_0_1_00_111_010_101_0_x_00;
      patterns[7939] = 33'b1000110101110010_1_1_00_111_010_101_0_x_00;
      patterns[7940] = 33'b1000110101110010_0_0_00_000_000_000_0_0_00;
      patterns[7941] = 33'b1001010101110010_0_1_01_111_010_101_0_x_00;
      patterns[7942] = 33'b1001110101110010_1_1_01_111_010_101_0_x_00;
      patterns[7943] = 33'b1001110101110010_0_0_00_000_000_000_0_0_00;
      patterns[7944] = 33'b1010010101110010_0_1_10_111_010_101_0_x_00;
      patterns[7945] = 33'b1010110101110010_1_1_10_111_010_101_0_x_00;
      patterns[7946] = 33'b1010110101110010_0_0_00_000_000_000_0_0_00;
      patterns[7947] = 33'b1011010101110010_0_1_11_111_010_101_0_x_00;
      patterns[7948] = 33'b1011110101110010_1_1_11_111_010_101_0_x_00;
      patterns[7949] = 33'b1011110101110010_0_0_00_000_000_000_0_0_00;
      patterns[7950] = 33'b0101010101110000_0_1_xx_111_xxx_101_0_1_01;
      patterns[7951] = 33'b0101110101110000_1_1_xx_111_xxx_101_0_1_01;
      patterns[7952] = 33'b0101110101110000_0_0_00_000_000_000_0_0_00;
      patterns[7953] = 33'b0100010101110000_0_0_xx_111_101_xxx_1_x_xx;
      patterns[7954] = 33'b0100110101110000_1_0_xx_111_101_xxx_1_x_xx;
      patterns[7955] = 33'b0100110101110000_0_0_00_000_000_000_0_0_00;
      patterns[7956] = 33'b0000010101000110_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7957] = 33'b0000110101000110_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7958] = 33'b0000110101000110_0_0_00_000_000_000_0_0_00;
      patterns[7959] = 33'b1000010101110011_0_1_00_111_011_101_0_x_00;
      patterns[7960] = 33'b1000110101110011_1_1_00_111_011_101_0_x_00;
      patterns[7961] = 33'b1000110101110011_0_0_00_000_000_000_0_0_00;
      patterns[7962] = 33'b1001010101110011_0_1_01_111_011_101_0_x_00;
      patterns[7963] = 33'b1001110101110011_1_1_01_111_011_101_0_x_00;
      patterns[7964] = 33'b1001110101110011_0_0_00_000_000_000_0_0_00;
      patterns[7965] = 33'b1010010101110011_0_1_10_111_011_101_0_x_00;
      patterns[7966] = 33'b1010110101110011_1_1_10_111_011_101_0_x_00;
      patterns[7967] = 33'b1010110101110011_0_0_00_000_000_000_0_0_00;
      patterns[7968] = 33'b1011010101110011_0_1_11_111_011_101_0_x_00;
      patterns[7969] = 33'b1011110101110011_1_1_11_111_011_101_0_x_00;
      patterns[7970] = 33'b1011110101110011_0_0_00_000_000_000_0_0_00;
      patterns[7971] = 33'b0101010101110000_0_1_xx_111_xxx_101_0_1_01;
      patterns[7972] = 33'b0101110101110000_1_1_xx_111_xxx_101_0_1_01;
      patterns[7973] = 33'b0101110101110000_0_0_00_000_000_000_0_0_00;
      patterns[7974] = 33'b0100010101110000_0_0_xx_111_101_xxx_1_x_xx;
      patterns[7975] = 33'b0100110101110000_1_0_xx_111_101_xxx_1_x_xx;
      patterns[7976] = 33'b0100110101110000_0_0_00_000_000_000_0_0_00;
      patterns[7977] = 33'b0000010111100010_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7978] = 33'b0000110111100010_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[7979] = 33'b0000110111100010_0_0_00_000_000_000_0_0_00;
      patterns[7980] = 33'b1000010101110100_0_1_00_111_100_101_0_x_00;
      patterns[7981] = 33'b1000110101110100_1_1_00_111_100_101_0_x_00;
      patterns[7982] = 33'b1000110101110100_0_0_00_000_000_000_0_0_00;
      patterns[7983] = 33'b1001010101110100_0_1_01_111_100_101_0_x_00;
      patterns[7984] = 33'b1001110101110100_1_1_01_111_100_101_0_x_00;
      patterns[7985] = 33'b1001110101110100_0_0_00_000_000_000_0_0_00;
      patterns[7986] = 33'b1010010101110100_0_1_10_111_100_101_0_x_00;
      patterns[7987] = 33'b1010110101110100_1_1_10_111_100_101_0_x_00;
      patterns[7988] = 33'b1010110101110100_0_0_00_000_000_000_0_0_00;
      patterns[7989] = 33'b1011010101110100_0_1_11_111_100_101_0_x_00;
      patterns[7990] = 33'b1011110101110100_1_1_11_111_100_101_0_x_00;
      patterns[7991] = 33'b1011110101110100_0_0_00_000_000_000_0_0_00;
      patterns[7992] = 33'b0101010101110000_0_1_xx_111_xxx_101_0_1_01;
      patterns[7993] = 33'b0101110101110000_1_1_xx_111_xxx_101_0_1_01;
      patterns[7994] = 33'b0101110101110000_0_0_00_000_000_000_0_0_00;
      patterns[7995] = 33'b0100010101110000_0_0_xx_111_101_xxx_1_x_xx;
      patterns[7996] = 33'b0100110101110000_1_0_xx_111_101_xxx_1_x_xx;
      patterns[7997] = 33'b0100110101110000_0_0_00_000_000_000_0_0_00;
      patterns[7998] = 33'b0000010101111100_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[7999] = 33'b0000110101111100_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[8000] = 33'b0000110101111100_0_0_00_000_000_000_0_0_00;
      patterns[8001] = 33'b1000010101110101_0_1_00_111_101_101_0_x_00;
      patterns[8002] = 33'b1000110101110101_1_1_00_111_101_101_0_x_00;
      patterns[8003] = 33'b1000110101110101_0_0_00_000_000_000_0_0_00;
      patterns[8004] = 33'b1001010101110101_0_1_01_111_101_101_0_x_00;
      patterns[8005] = 33'b1001110101110101_1_1_01_111_101_101_0_x_00;
      patterns[8006] = 33'b1001110101110101_0_0_00_000_000_000_0_0_00;
      patterns[8007] = 33'b1010010101110101_0_1_10_111_101_101_0_x_00;
      patterns[8008] = 33'b1010110101110101_1_1_10_111_101_101_0_x_00;
      patterns[8009] = 33'b1010110101110101_0_0_00_000_000_000_0_0_00;
      patterns[8010] = 33'b1011010101110101_0_1_11_111_101_101_0_x_00;
      patterns[8011] = 33'b1011110101110101_1_1_11_111_101_101_0_x_00;
      patterns[8012] = 33'b1011110101110101_0_0_00_000_000_000_0_0_00;
      patterns[8013] = 33'b0101010101110000_0_1_xx_111_xxx_101_0_1_01;
      patterns[8014] = 33'b0101110101110000_1_1_xx_111_xxx_101_0_1_01;
      patterns[8015] = 33'b0101110101110000_0_0_00_000_000_000_0_0_00;
      patterns[8016] = 33'b0100010101110000_0_0_xx_111_101_xxx_1_x_xx;
      patterns[8017] = 33'b0100110101110000_1_0_xx_111_101_xxx_1_x_xx;
      patterns[8018] = 33'b0100110101110000_0_0_00_000_000_000_0_0_00;
      patterns[8019] = 33'b0000010111010010_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[8020] = 33'b0000110111010010_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[8021] = 33'b0000110111010010_0_0_00_000_000_000_0_0_00;
      patterns[8022] = 33'b1000010101110110_0_1_00_111_110_101_0_x_00;
      patterns[8023] = 33'b1000110101110110_1_1_00_111_110_101_0_x_00;
      patterns[8024] = 33'b1000110101110110_0_0_00_000_000_000_0_0_00;
      patterns[8025] = 33'b1001010101110110_0_1_01_111_110_101_0_x_00;
      patterns[8026] = 33'b1001110101110110_1_1_01_111_110_101_0_x_00;
      patterns[8027] = 33'b1001110101110110_0_0_00_000_000_000_0_0_00;
      patterns[8028] = 33'b1010010101110110_0_1_10_111_110_101_0_x_00;
      patterns[8029] = 33'b1010110101110110_1_1_10_111_110_101_0_x_00;
      patterns[8030] = 33'b1010110101110110_0_0_00_000_000_000_0_0_00;
      patterns[8031] = 33'b1011010101110110_0_1_11_111_110_101_0_x_00;
      patterns[8032] = 33'b1011110101110110_1_1_11_111_110_101_0_x_00;
      patterns[8033] = 33'b1011110101110110_0_0_00_000_000_000_0_0_00;
      patterns[8034] = 33'b0101010101110000_0_1_xx_111_xxx_101_0_1_01;
      patterns[8035] = 33'b0101110101110000_1_1_xx_111_xxx_101_0_1_01;
      patterns[8036] = 33'b0101110101110000_0_0_00_000_000_000_0_0_00;
      patterns[8037] = 33'b0100010101110000_0_0_xx_111_101_xxx_1_x_xx;
      patterns[8038] = 33'b0100110101110000_1_0_xx_111_101_xxx_1_x_xx;
      patterns[8039] = 33'b0100110101110000_0_0_00_000_000_000_0_0_00;
      patterns[8040] = 33'b0000010111010001_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[8041] = 33'b0000110111010001_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[8042] = 33'b0000110111010001_0_0_00_000_000_000_0_0_00;
      patterns[8043] = 33'b1000010101110111_0_1_00_111_111_101_0_x_00;
      patterns[8044] = 33'b1000110101110111_1_1_00_111_111_101_0_x_00;
      patterns[8045] = 33'b1000110101110111_0_0_00_000_000_000_0_0_00;
      patterns[8046] = 33'b1001010101110111_0_1_01_111_111_101_0_x_00;
      patterns[8047] = 33'b1001110101110111_1_1_01_111_111_101_0_x_00;
      patterns[8048] = 33'b1001110101110111_0_0_00_000_000_000_0_0_00;
      patterns[8049] = 33'b1010010101110111_0_1_10_111_111_101_0_x_00;
      patterns[8050] = 33'b1010110101110111_1_1_10_111_111_101_0_x_00;
      patterns[8051] = 33'b1010110101110111_0_0_00_000_000_000_0_0_00;
      patterns[8052] = 33'b1011010101110111_0_1_11_111_111_101_0_x_00;
      patterns[8053] = 33'b1011110101110111_1_1_11_111_111_101_0_x_00;
      patterns[8054] = 33'b1011110101110111_0_0_00_000_000_000_0_0_00;
      patterns[8055] = 33'b0101010101110000_0_1_xx_111_xxx_101_0_1_01;
      patterns[8056] = 33'b0101110101110000_1_1_xx_111_xxx_101_0_1_01;
      patterns[8057] = 33'b0101110101110000_0_0_00_000_000_000_0_0_00;
      patterns[8058] = 33'b0100010101110000_0_0_xx_111_101_xxx_1_x_xx;
      patterns[8059] = 33'b0100110101110000_1_0_xx_111_101_xxx_1_x_xx;
      patterns[8060] = 33'b0100110101110000_0_0_00_000_000_000_0_0_00;
      patterns[8061] = 33'b0000010100000010_0_1_xx_xxx_xxx_101_0_x_10;
      patterns[8062] = 33'b0000110100000010_1_1_xx_xxx_xxx_101_0_x_10;
      patterns[8063] = 33'b0000110100000010_0_0_00_000_000_000_0_0_00;
      patterns[8064] = 33'b1000011000000000_0_1_00_000_000_110_0_x_00;
      patterns[8065] = 33'b1000111000000000_1_1_00_000_000_110_0_x_00;
      patterns[8066] = 33'b1000111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8067] = 33'b1001011000000000_0_1_01_000_000_110_0_x_00;
      patterns[8068] = 33'b1001111000000000_1_1_01_000_000_110_0_x_00;
      patterns[8069] = 33'b1001111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8070] = 33'b1010011000000000_0_1_10_000_000_110_0_x_00;
      patterns[8071] = 33'b1010111000000000_1_1_10_000_000_110_0_x_00;
      patterns[8072] = 33'b1010111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8073] = 33'b1011011000000000_0_1_11_000_000_110_0_x_00;
      patterns[8074] = 33'b1011111000000000_1_1_11_000_000_110_0_x_00;
      patterns[8075] = 33'b1011111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8076] = 33'b0101011000000000_0_1_xx_000_xxx_110_0_1_01;
      patterns[8077] = 33'b0101111000000000_1_1_xx_000_xxx_110_0_1_01;
      patterns[8078] = 33'b0101111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8079] = 33'b0100011000000000_0_0_xx_000_110_xxx_1_x_xx;
      patterns[8080] = 33'b0100111000000000_1_0_xx_000_110_xxx_1_x_xx;
      patterns[8081] = 33'b0100111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8082] = 33'b0000011011011011_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8083] = 33'b0000111011011011_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8084] = 33'b0000111011011011_0_0_00_000_000_000_0_0_00;
      patterns[8085] = 33'b1000011000000001_0_1_00_000_001_110_0_x_00;
      patterns[8086] = 33'b1000111000000001_1_1_00_000_001_110_0_x_00;
      patterns[8087] = 33'b1000111000000001_0_0_00_000_000_000_0_0_00;
      patterns[8088] = 33'b1001011000000001_0_1_01_000_001_110_0_x_00;
      patterns[8089] = 33'b1001111000000001_1_1_01_000_001_110_0_x_00;
      patterns[8090] = 33'b1001111000000001_0_0_00_000_000_000_0_0_00;
      patterns[8091] = 33'b1010011000000001_0_1_10_000_001_110_0_x_00;
      patterns[8092] = 33'b1010111000000001_1_1_10_000_001_110_0_x_00;
      patterns[8093] = 33'b1010111000000001_0_0_00_000_000_000_0_0_00;
      patterns[8094] = 33'b1011011000000001_0_1_11_000_001_110_0_x_00;
      patterns[8095] = 33'b1011111000000001_1_1_11_000_001_110_0_x_00;
      patterns[8096] = 33'b1011111000000001_0_0_00_000_000_000_0_0_00;
      patterns[8097] = 33'b0101011000000000_0_1_xx_000_xxx_110_0_1_01;
      patterns[8098] = 33'b0101111000000000_1_1_xx_000_xxx_110_0_1_01;
      patterns[8099] = 33'b0101111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8100] = 33'b0100011000000000_0_0_xx_000_110_xxx_1_x_xx;
      patterns[8101] = 33'b0100111000000000_1_0_xx_000_110_xxx_1_x_xx;
      patterns[8102] = 33'b0100111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8103] = 33'b0000011010110110_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8104] = 33'b0000111010110110_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8105] = 33'b0000111010110110_0_0_00_000_000_000_0_0_00;
      patterns[8106] = 33'b1000011000000010_0_1_00_000_010_110_0_x_00;
      patterns[8107] = 33'b1000111000000010_1_1_00_000_010_110_0_x_00;
      patterns[8108] = 33'b1000111000000010_0_0_00_000_000_000_0_0_00;
      patterns[8109] = 33'b1001011000000010_0_1_01_000_010_110_0_x_00;
      patterns[8110] = 33'b1001111000000010_1_1_01_000_010_110_0_x_00;
      patterns[8111] = 33'b1001111000000010_0_0_00_000_000_000_0_0_00;
      patterns[8112] = 33'b1010011000000010_0_1_10_000_010_110_0_x_00;
      patterns[8113] = 33'b1010111000000010_1_1_10_000_010_110_0_x_00;
      patterns[8114] = 33'b1010111000000010_0_0_00_000_000_000_0_0_00;
      patterns[8115] = 33'b1011011000000010_0_1_11_000_010_110_0_x_00;
      patterns[8116] = 33'b1011111000000010_1_1_11_000_010_110_0_x_00;
      patterns[8117] = 33'b1011111000000010_0_0_00_000_000_000_0_0_00;
      patterns[8118] = 33'b0101011000000000_0_1_xx_000_xxx_110_0_1_01;
      patterns[8119] = 33'b0101111000000000_1_1_xx_000_xxx_110_0_1_01;
      patterns[8120] = 33'b0101111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8121] = 33'b0100011000000000_0_0_xx_000_110_xxx_1_x_xx;
      patterns[8122] = 33'b0100111000000000_1_0_xx_000_110_xxx_1_x_xx;
      patterns[8123] = 33'b0100111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8124] = 33'b0000011011100110_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8125] = 33'b0000111011100110_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8126] = 33'b0000111011100110_0_0_00_000_000_000_0_0_00;
      patterns[8127] = 33'b1000011000000011_0_1_00_000_011_110_0_x_00;
      patterns[8128] = 33'b1000111000000011_1_1_00_000_011_110_0_x_00;
      patterns[8129] = 33'b1000111000000011_0_0_00_000_000_000_0_0_00;
      patterns[8130] = 33'b1001011000000011_0_1_01_000_011_110_0_x_00;
      patterns[8131] = 33'b1001111000000011_1_1_01_000_011_110_0_x_00;
      patterns[8132] = 33'b1001111000000011_0_0_00_000_000_000_0_0_00;
      patterns[8133] = 33'b1010011000000011_0_1_10_000_011_110_0_x_00;
      patterns[8134] = 33'b1010111000000011_1_1_10_000_011_110_0_x_00;
      patterns[8135] = 33'b1010111000000011_0_0_00_000_000_000_0_0_00;
      patterns[8136] = 33'b1011011000000011_0_1_11_000_011_110_0_x_00;
      patterns[8137] = 33'b1011111000000011_1_1_11_000_011_110_0_x_00;
      patterns[8138] = 33'b1011111000000011_0_0_00_000_000_000_0_0_00;
      patterns[8139] = 33'b0101011000000000_0_1_xx_000_xxx_110_0_1_01;
      patterns[8140] = 33'b0101111000000000_1_1_xx_000_xxx_110_0_1_01;
      patterns[8141] = 33'b0101111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8142] = 33'b0100011000000000_0_0_xx_000_110_xxx_1_x_xx;
      patterns[8143] = 33'b0100111000000000_1_0_xx_000_110_xxx_1_x_xx;
      patterns[8144] = 33'b0100111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8145] = 33'b0000011010001000_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8146] = 33'b0000111010001000_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8147] = 33'b0000111010001000_0_0_00_000_000_000_0_0_00;
      patterns[8148] = 33'b1000011000000100_0_1_00_000_100_110_0_x_00;
      patterns[8149] = 33'b1000111000000100_1_1_00_000_100_110_0_x_00;
      patterns[8150] = 33'b1000111000000100_0_0_00_000_000_000_0_0_00;
      patterns[8151] = 33'b1001011000000100_0_1_01_000_100_110_0_x_00;
      patterns[8152] = 33'b1001111000000100_1_1_01_000_100_110_0_x_00;
      patterns[8153] = 33'b1001111000000100_0_0_00_000_000_000_0_0_00;
      patterns[8154] = 33'b1010011000000100_0_1_10_000_100_110_0_x_00;
      patterns[8155] = 33'b1010111000000100_1_1_10_000_100_110_0_x_00;
      patterns[8156] = 33'b1010111000000100_0_0_00_000_000_000_0_0_00;
      patterns[8157] = 33'b1011011000000100_0_1_11_000_100_110_0_x_00;
      patterns[8158] = 33'b1011111000000100_1_1_11_000_100_110_0_x_00;
      patterns[8159] = 33'b1011111000000100_0_0_00_000_000_000_0_0_00;
      patterns[8160] = 33'b0101011000000000_0_1_xx_000_xxx_110_0_1_01;
      patterns[8161] = 33'b0101111000000000_1_1_xx_000_xxx_110_0_1_01;
      patterns[8162] = 33'b0101111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8163] = 33'b0100011000000000_0_0_xx_000_110_xxx_1_x_xx;
      patterns[8164] = 33'b0100111000000000_1_0_xx_000_110_xxx_1_x_xx;
      patterns[8165] = 33'b0100111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8166] = 33'b0000011001000100_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8167] = 33'b0000111001000100_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8168] = 33'b0000111001000100_0_0_00_000_000_000_0_0_00;
      patterns[8169] = 33'b1000011000000101_0_1_00_000_101_110_0_x_00;
      patterns[8170] = 33'b1000111000000101_1_1_00_000_101_110_0_x_00;
      patterns[8171] = 33'b1000111000000101_0_0_00_000_000_000_0_0_00;
      patterns[8172] = 33'b1001011000000101_0_1_01_000_101_110_0_x_00;
      patterns[8173] = 33'b1001111000000101_1_1_01_000_101_110_0_x_00;
      patterns[8174] = 33'b1001111000000101_0_0_00_000_000_000_0_0_00;
      patterns[8175] = 33'b1010011000000101_0_1_10_000_101_110_0_x_00;
      patterns[8176] = 33'b1010111000000101_1_1_10_000_101_110_0_x_00;
      patterns[8177] = 33'b1010111000000101_0_0_00_000_000_000_0_0_00;
      patterns[8178] = 33'b1011011000000101_0_1_11_000_101_110_0_x_00;
      patterns[8179] = 33'b1011111000000101_1_1_11_000_101_110_0_x_00;
      patterns[8180] = 33'b1011111000000101_0_0_00_000_000_000_0_0_00;
      patterns[8181] = 33'b0101011000000000_0_1_xx_000_xxx_110_0_1_01;
      patterns[8182] = 33'b0101111000000000_1_1_xx_000_xxx_110_0_1_01;
      patterns[8183] = 33'b0101111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8184] = 33'b0100011000000000_0_0_xx_000_110_xxx_1_x_xx;
      patterns[8185] = 33'b0100111000000000_1_0_xx_000_110_xxx_1_x_xx;
      patterns[8186] = 33'b0100111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8187] = 33'b0000011001101100_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8188] = 33'b0000111001101100_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8189] = 33'b0000111001101100_0_0_00_000_000_000_0_0_00;
      patterns[8190] = 33'b1000011000000110_0_1_00_000_110_110_0_x_00;
      patterns[8191] = 33'b1000111000000110_1_1_00_000_110_110_0_x_00;
      patterns[8192] = 33'b1000111000000110_0_0_00_000_000_000_0_0_00;
      patterns[8193] = 33'b1001011000000110_0_1_01_000_110_110_0_x_00;
      patterns[8194] = 33'b1001111000000110_1_1_01_000_110_110_0_x_00;
      patterns[8195] = 33'b1001111000000110_0_0_00_000_000_000_0_0_00;
      patterns[8196] = 33'b1010011000000110_0_1_10_000_110_110_0_x_00;
      patterns[8197] = 33'b1010111000000110_1_1_10_000_110_110_0_x_00;
      patterns[8198] = 33'b1010111000000110_0_0_00_000_000_000_0_0_00;
      patterns[8199] = 33'b1011011000000110_0_1_11_000_110_110_0_x_00;
      patterns[8200] = 33'b1011111000000110_1_1_11_000_110_110_0_x_00;
      patterns[8201] = 33'b1011111000000110_0_0_00_000_000_000_0_0_00;
      patterns[8202] = 33'b0101011000000000_0_1_xx_000_xxx_110_0_1_01;
      patterns[8203] = 33'b0101111000000000_1_1_xx_000_xxx_110_0_1_01;
      patterns[8204] = 33'b0101111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8205] = 33'b0100011000000000_0_0_xx_000_110_xxx_1_x_xx;
      patterns[8206] = 33'b0100111000000000_1_0_xx_000_110_xxx_1_x_xx;
      patterns[8207] = 33'b0100111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8208] = 33'b0000011011011111_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8209] = 33'b0000111011011111_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8210] = 33'b0000111011011111_0_0_00_000_000_000_0_0_00;
      patterns[8211] = 33'b1000011000000111_0_1_00_000_111_110_0_x_00;
      patterns[8212] = 33'b1000111000000111_1_1_00_000_111_110_0_x_00;
      patterns[8213] = 33'b1000111000000111_0_0_00_000_000_000_0_0_00;
      patterns[8214] = 33'b1001011000000111_0_1_01_000_111_110_0_x_00;
      patterns[8215] = 33'b1001111000000111_1_1_01_000_111_110_0_x_00;
      patterns[8216] = 33'b1001111000000111_0_0_00_000_000_000_0_0_00;
      patterns[8217] = 33'b1010011000000111_0_1_10_000_111_110_0_x_00;
      patterns[8218] = 33'b1010111000000111_1_1_10_000_111_110_0_x_00;
      patterns[8219] = 33'b1010111000000111_0_0_00_000_000_000_0_0_00;
      patterns[8220] = 33'b1011011000000111_0_1_11_000_111_110_0_x_00;
      patterns[8221] = 33'b1011111000000111_1_1_11_000_111_110_0_x_00;
      patterns[8222] = 33'b1011111000000111_0_0_00_000_000_000_0_0_00;
      patterns[8223] = 33'b0101011000000000_0_1_xx_000_xxx_110_0_1_01;
      patterns[8224] = 33'b0101111000000000_1_1_xx_000_xxx_110_0_1_01;
      patterns[8225] = 33'b0101111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8226] = 33'b0100011000000000_0_0_xx_000_110_xxx_1_x_xx;
      patterns[8227] = 33'b0100111000000000_1_0_xx_000_110_xxx_1_x_xx;
      patterns[8228] = 33'b0100111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8229] = 33'b0000011001000001_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8230] = 33'b0000111001000001_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8231] = 33'b0000111001000001_0_0_00_000_000_000_0_0_00;
      patterns[8232] = 33'b1000011000010000_0_1_00_001_000_110_0_x_00;
      patterns[8233] = 33'b1000111000010000_1_1_00_001_000_110_0_x_00;
      patterns[8234] = 33'b1000111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8235] = 33'b1001011000010000_0_1_01_001_000_110_0_x_00;
      patterns[8236] = 33'b1001111000010000_1_1_01_001_000_110_0_x_00;
      patterns[8237] = 33'b1001111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8238] = 33'b1010011000010000_0_1_10_001_000_110_0_x_00;
      patterns[8239] = 33'b1010111000010000_1_1_10_001_000_110_0_x_00;
      patterns[8240] = 33'b1010111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8241] = 33'b1011011000010000_0_1_11_001_000_110_0_x_00;
      patterns[8242] = 33'b1011111000010000_1_1_11_001_000_110_0_x_00;
      patterns[8243] = 33'b1011111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8244] = 33'b0101011000010000_0_1_xx_001_xxx_110_0_1_01;
      patterns[8245] = 33'b0101111000010000_1_1_xx_001_xxx_110_0_1_01;
      patterns[8246] = 33'b0101111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8247] = 33'b0100011000010000_0_0_xx_001_110_xxx_1_x_xx;
      patterns[8248] = 33'b0100111000010000_1_0_xx_001_110_xxx_1_x_xx;
      patterns[8249] = 33'b0100111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8250] = 33'b0000011011110001_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8251] = 33'b0000111011110001_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8252] = 33'b0000111011110001_0_0_00_000_000_000_0_0_00;
      patterns[8253] = 33'b1000011000010001_0_1_00_001_001_110_0_x_00;
      patterns[8254] = 33'b1000111000010001_1_1_00_001_001_110_0_x_00;
      patterns[8255] = 33'b1000111000010001_0_0_00_000_000_000_0_0_00;
      patterns[8256] = 33'b1001011000010001_0_1_01_001_001_110_0_x_00;
      patterns[8257] = 33'b1001111000010001_1_1_01_001_001_110_0_x_00;
      patterns[8258] = 33'b1001111000010001_0_0_00_000_000_000_0_0_00;
      patterns[8259] = 33'b1010011000010001_0_1_10_001_001_110_0_x_00;
      patterns[8260] = 33'b1010111000010001_1_1_10_001_001_110_0_x_00;
      patterns[8261] = 33'b1010111000010001_0_0_00_000_000_000_0_0_00;
      patterns[8262] = 33'b1011011000010001_0_1_11_001_001_110_0_x_00;
      patterns[8263] = 33'b1011111000010001_1_1_11_001_001_110_0_x_00;
      patterns[8264] = 33'b1011111000010001_0_0_00_000_000_000_0_0_00;
      patterns[8265] = 33'b0101011000010000_0_1_xx_001_xxx_110_0_1_01;
      patterns[8266] = 33'b0101111000010000_1_1_xx_001_xxx_110_0_1_01;
      patterns[8267] = 33'b0101111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8268] = 33'b0100011000010000_0_0_xx_001_110_xxx_1_x_xx;
      patterns[8269] = 33'b0100111000010000_1_0_xx_001_110_xxx_1_x_xx;
      patterns[8270] = 33'b0100111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8271] = 33'b0000011001001111_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8272] = 33'b0000111001001111_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8273] = 33'b0000111001001111_0_0_00_000_000_000_0_0_00;
      patterns[8274] = 33'b1000011000010010_0_1_00_001_010_110_0_x_00;
      patterns[8275] = 33'b1000111000010010_1_1_00_001_010_110_0_x_00;
      patterns[8276] = 33'b1000111000010010_0_0_00_000_000_000_0_0_00;
      patterns[8277] = 33'b1001011000010010_0_1_01_001_010_110_0_x_00;
      patterns[8278] = 33'b1001111000010010_1_1_01_001_010_110_0_x_00;
      patterns[8279] = 33'b1001111000010010_0_0_00_000_000_000_0_0_00;
      patterns[8280] = 33'b1010011000010010_0_1_10_001_010_110_0_x_00;
      patterns[8281] = 33'b1010111000010010_1_1_10_001_010_110_0_x_00;
      patterns[8282] = 33'b1010111000010010_0_0_00_000_000_000_0_0_00;
      patterns[8283] = 33'b1011011000010010_0_1_11_001_010_110_0_x_00;
      patterns[8284] = 33'b1011111000010010_1_1_11_001_010_110_0_x_00;
      patterns[8285] = 33'b1011111000010010_0_0_00_000_000_000_0_0_00;
      patterns[8286] = 33'b0101011000010000_0_1_xx_001_xxx_110_0_1_01;
      patterns[8287] = 33'b0101111000010000_1_1_xx_001_xxx_110_0_1_01;
      patterns[8288] = 33'b0101111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8289] = 33'b0100011000010000_0_0_xx_001_110_xxx_1_x_xx;
      patterns[8290] = 33'b0100111000010000_1_0_xx_001_110_xxx_1_x_xx;
      patterns[8291] = 33'b0100111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8292] = 33'b0000011000001010_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8293] = 33'b0000111000001010_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8294] = 33'b0000111000001010_0_0_00_000_000_000_0_0_00;
      patterns[8295] = 33'b1000011000010011_0_1_00_001_011_110_0_x_00;
      patterns[8296] = 33'b1000111000010011_1_1_00_001_011_110_0_x_00;
      patterns[8297] = 33'b1000111000010011_0_0_00_000_000_000_0_0_00;
      patterns[8298] = 33'b1001011000010011_0_1_01_001_011_110_0_x_00;
      patterns[8299] = 33'b1001111000010011_1_1_01_001_011_110_0_x_00;
      patterns[8300] = 33'b1001111000010011_0_0_00_000_000_000_0_0_00;
      patterns[8301] = 33'b1010011000010011_0_1_10_001_011_110_0_x_00;
      patterns[8302] = 33'b1010111000010011_1_1_10_001_011_110_0_x_00;
      patterns[8303] = 33'b1010111000010011_0_0_00_000_000_000_0_0_00;
      patterns[8304] = 33'b1011011000010011_0_1_11_001_011_110_0_x_00;
      patterns[8305] = 33'b1011111000010011_1_1_11_001_011_110_0_x_00;
      patterns[8306] = 33'b1011111000010011_0_0_00_000_000_000_0_0_00;
      patterns[8307] = 33'b0101011000010000_0_1_xx_001_xxx_110_0_1_01;
      patterns[8308] = 33'b0101111000010000_1_1_xx_001_xxx_110_0_1_01;
      patterns[8309] = 33'b0101111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8310] = 33'b0100011000010000_0_0_xx_001_110_xxx_1_x_xx;
      patterns[8311] = 33'b0100111000010000_1_0_xx_001_110_xxx_1_x_xx;
      patterns[8312] = 33'b0100111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8313] = 33'b0000011011111000_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8314] = 33'b0000111011111000_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8315] = 33'b0000111011111000_0_0_00_000_000_000_0_0_00;
      patterns[8316] = 33'b1000011000010100_0_1_00_001_100_110_0_x_00;
      patterns[8317] = 33'b1000111000010100_1_1_00_001_100_110_0_x_00;
      patterns[8318] = 33'b1000111000010100_0_0_00_000_000_000_0_0_00;
      patterns[8319] = 33'b1001011000010100_0_1_01_001_100_110_0_x_00;
      patterns[8320] = 33'b1001111000010100_1_1_01_001_100_110_0_x_00;
      patterns[8321] = 33'b1001111000010100_0_0_00_000_000_000_0_0_00;
      patterns[8322] = 33'b1010011000010100_0_1_10_001_100_110_0_x_00;
      patterns[8323] = 33'b1010111000010100_1_1_10_001_100_110_0_x_00;
      patterns[8324] = 33'b1010111000010100_0_0_00_000_000_000_0_0_00;
      patterns[8325] = 33'b1011011000010100_0_1_11_001_100_110_0_x_00;
      patterns[8326] = 33'b1011111000010100_1_1_11_001_100_110_0_x_00;
      patterns[8327] = 33'b1011111000010100_0_0_00_000_000_000_0_0_00;
      patterns[8328] = 33'b0101011000010000_0_1_xx_001_xxx_110_0_1_01;
      patterns[8329] = 33'b0101111000010000_1_1_xx_001_xxx_110_0_1_01;
      patterns[8330] = 33'b0101111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8331] = 33'b0100011000010000_0_0_xx_001_110_xxx_1_x_xx;
      patterns[8332] = 33'b0100111000010000_1_0_xx_001_110_xxx_1_x_xx;
      patterns[8333] = 33'b0100111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8334] = 33'b0000011000000000_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8335] = 33'b0000111000000000_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8336] = 33'b0000111000000000_0_0_00_000_000_000_0_0_00;
      patterns[8337] = 33'b1000011000010101_0_1_00_001_101_110_0_x_00;
      patterns[8338] = 33'b1000111000010101_1_1_00_001_101_110_0_x_00;
      patterns[8339] = 33'b1000111000010101_0_0_00_000_000_000_0_0_00;
      patterns[8340] = 33'b1001011000010101_0_1_01_001_101_110_0_x_00;
      patterns[8341] = 33'b1001111000010101_1_1_01_001_101_110_0_x_00;
      patterns[8342] = 33'b1001111000010101_0_0_00_000_000_000_0_0_00;
      patterns[8343] = 33'b1010011000010101_0_1_10_001_101_110_0_x_00;
      patterns[8344] = 33'b1010111000010101_1_1_10_001_101_110_0_x_00;
      patterns[8345] = 33'b1010111000010101_0_0_00_000_000_000_0_0_00;
      patterns[8346] = 33'b1011011000010101_0_1_11_001_101_110_0_x_00;
      patterns[8347] = 33'b1011111000010101_1_1_11_001_101_110_0_x_00;
      patterns[8348] = 33'b1011111000010101_0_0_00_000_000_000_0_0_00;
      patterns[8349] = 33'b0101011000010000_0_1_xx_001_xxx_110_0_1_01;
      patterns[8350] = 33'b0101111000010000_1_1_xx_001_xxx_110_0_1_01;
      patterns[8351] = 33'b0101111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8352] = 33'b0100011000010000_0_0_xx_001_110_xxx_1_x_xx;
      patterns[8353] = 33'b0100111000010000_1_0_xx_001_110_xxx_1_x_xx;
      patterns[8354] = 33'b0100111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8355] = 33'b0000011011010010_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8356] = 33'b0000111011010010_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8357] = 33'b0000111011010010_0_0_00_000_000_000_0_0_00;
      patterns[8358] = 33'b1000011000010110_0_1_00_001_110_110_0_x_00;
      patterns[8359] = 33'b1000111000010110_1_1_00_001_110_110_0_x_00;
      patterns[8360] = 33'b1000111000010110_0_0_00_000_000_000_0_0_00;
      patterns[8361] = 33'b1001011000010110_0_1_01_001_110_110_0_x_00;
      patterns[8362] = 33'b1001111000010110_1_1_01_001_110_110_0_x_00;
      patterns[8363] = 33'b1001111000010110_0_0_00_000_000_000_0_0_00;
      patterns[8364] = 33'b1010011000010110_0_1_10_001_110_110_0_x_00;
      patterns[8365] = 33'b1010111000010110_1_1_10_001_110_110_0_x_00;
      patterns[8366] = 33'b1010111000010110_0_0_00_000_000_000_0_0_00;
      patterns[8367] = 33'b1011011000010110_0_1_11_001_110_110_0_x_00;
      patterns[8368] = 33'b1011111000010110_1_1_11_001_110_110_0_x_00;
      patterns[8369] = 33'b1011111000010110_0_0_00_000_000_000_0_0_00;
      patterns[8370] = 33'b0101011000010000_0_1_xx_001_xxx_110_0_1_01;
      patterns[8371] = 33'b0101111000010000_1_1_xx_001_xxx_110_0_1_01;
      patterns[8372] = 33'b0101111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8373] = 33'b0100011000010000_0_0_xx_001_110_xxx_1_x_xx;
      patterns[8374] = 33'b0100111000010000_1_0_xx_001_110_xxx_1_x_xx;
      patterns[8375] = 33'b0100111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8376] = 33'b0000011000001001_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8377] = 33'b0000111000001001_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8378] = 33'b0000111000001001_0_0_00_000_000_000_0_0_00;
      patterns[8379] = 33'b1000011000010111_0_1_00_001_111_110_0_x_00;
      patterns[8380] = 33'b1000111000010111_1_1_00_001_111_110_0_x_00;
      patterns[8381] = 33'b1000111000010111_0_0_00_000_000_000_0_0_00;
      patterns[8382] = 33'b1001011000010111_0_1_01_001_111_110_0_x_00;
      patterns[8383] = 33'b1001111000010111_1_1_01_001_111_110_0_x_00;
      patterns[8384] = 33'b1001111000010111_0_0_00_000_000_000_0_0_00;
      patterns[8385] = 33'b1010011000010111_0_1_10_001_111_110_0_x_00;
      patterns[8386] = 33'b1010111000010111_1_1_10_001_111_110_0_x_00;
      patterns[8387] = 33'b1010111000010111_0_0_00_000_000_000_0_0_00;
      patterns[8388] = 33'b1011011000010111_0_1_11_001_111_110_0_x_00;
      patterns[8389] = 33'b1011111000010111_1_1_11_001_111_110_0_x_00;
      patterns[8390] = 33'b1011111000010111_0_0_00_000_000_000_0_0_00;
      patterns[8391] = 33'b0101011000010000_0_1_xx_001_xxx_110_0_1_01;
      patterns[8392] = 33'b0101111000010000_1_1_xx_001_xxx_110_0_1_01;
      patterns[8393] = 33'b0101111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8394] = 33'b0100011000010000_0_0_xx_001_110_xxx_1_x_xx;
      patterns[8395] = 33'b0100111000010000_1_0_xx_001_110_xxx_1_x_xx;
      patterns[8396] = 33'b0100111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8397] = 33'b0000011000101110_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8398] = 33'b0000111000101110_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8399] = 33'b0000111000101110_0_0_00_000_000_000_0_0_00;
      patterns[8400] = 33'b1000011000100000_0_1_00_010_000_110_0_x_00;
      patterns[8401] = 33'b1000111000100000_1_1_00_010_000_110_0_x_00;
      patterns[8402] = 33'b1000111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8403] = 33'b1001011000100000_0_1_01_010_000_110_0_x_00;
      patterns[8404] = 33'b1001111000100000_1_1_01_010_000_110_0_x_00;
      patterns[8405] = 33'b1001111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8406] = 33'b1010011000100000_0_1_10_010_000_110_0_x_00;
      patterns[8407] = 33'b1010111000100000_1_1_10_010_000_110_0_x_00;
      patterns[8408] = 33'b1010111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8409] = 33'b1011011000100000_0_1_11_010_000_110_0_x_00;
      patterns[8410] = 33'b1011111000100000_1_1_11_010_000_110_0_x_00;
      patterns[8411] = 33'b1011111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8412] = 33'b0101011000100000_0_1_xx_010_xxx_110_0_1_01;
      patterns[8413] = 33'b0101111000100000_1_1_xx_010_xxx_110_0_1_01;
      patterns[8414] = 33'b0101111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8415] = 33'b0100011000100000_0_0_xx_010_110_xxx_1_x_xx;
      patterns[8416] = 33'b0100111000100000_1_0_xx_010_110_xxx_1_x_xx;
      patterns[8417] = 33'b0100111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8418] = 33'b0000011000110110_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8419] = 33'b0000111000110110_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8420] = 33'b0000111000110110_0_0_00_000_000_000_0_0_00;
      patterns[8421] = 33'b1000011000100001_0_1_00_010_001_110_0_x_00;
      patterns[8422] = 33'b1000111000100001_1_1_00_010_001_110_0_x_00;
      patterns[8423] = 33'b1000111000100001_0_0_00_000_000_000_0_0_00;
      patterns[8424] = 33'b1001011000100001_0_1_01_010_001_110_0_x_00;
      patterns[8425] = 33'b1001111000100001_1_1_01_010_001_110_0_x_00;
      patterns[8426] = 33'b1001111000100001_0_0_00_000_000_000_0_0_00;
      patterns[8427] = 33'b1010011000100001_0_1_10_010_001_110_0_x_00;
      patterns[8428] = 33'b1010111000100001_1_1_10_010_001_110_0_x_00;
      patterns[8429] = 33'b1010111000100001_0_0_00_000_000_000_0_0_00;
      patterns[8430] = 33'b1011011000100001_0_1_11_010_001_110_0_x_00;
      patterns[8431] = 33'b1011111000100001_1_1_11_010_001_110_0_x_00;
      patterns[8432] = 33'b1011111000100001_0_0_00_000_000_000_0_0_00;
      patterns[8433] = 33'b0101011000100000_0_1_xx_010_xxx_110_0_1_01;
      patterns[8434] = 33'b0101111000100000_1_1_xx_010_xxx_110_0_1_01;
      patterns[8435] = 33'b0101111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8436] = 33'b0100011000100000_0_0_xx_010_110_xxx_1_x_xx;
      patterns[8437] = 33'b0100111000100000_1_0_xx_010_110_xxx_1_x_xx;
      patterns[8438] = 33'b0100111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8439] = 33'b0000011001001101_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8440] = 33'b0000111001001101_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8441] = 33'b0000111001001101_0_0_00_000_000_000_0_0_00;
      patterns[8442] = 33'b1000011000100010_0_1_00_010_010_110_0_x_00;
      patterns[8443] = 33'b1000111000100010_1_1_00_010_010_110_0_x_00;
      patterns[8444] = 33'b1000111000100010_0_0_00_000_000_000_0_0_00;
      patterns[8445] = 33'b1001011000100010_0_1_01_010_010_110_0_x_00;
      patterns[8446] = 33'b1001111000100010_1_1_01_010_010_110_0_x_00;
      patterns[8447] = 33'b1001111000100010_0_0_00_000_000_000_0_0_00;
      patterns[8448] = 33'b1010011000100010_0_1_10_010_010_110_0_x_00;
      patterns[8449] = 33'b1010111000100010_1_1_10_010_010_110_0_x_00;
      patterns[8450] = 33'b1010111000100010_0_0_00_000_000_000_0_0_00;
      patterns[8451] = 33'b1011011000100010_0_1_11_010_010_110_0_x_00;
      patterns[8452] = 33'b1011111000100010_1_1_11_010_010_110_0_x_00;
      patterns[8453] = 33'b1011111000100010_0_0_00_000_000_000_0_0_00;
      patterns[8454] = 33'b0101011000100000_0_1_xx_010_xxx_110_0_1_01;
      patterns[8455] = 33'b0101111000100000_1_1_xx_010_xxx_110_0_1_01;
      patterns[8456] = 33'b0101111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8457] = 33'b0100011000100000_0_0_xx_010_110_xxx_1_x_xx;
      patterns[8458] = 33'b0100111000100000_1_0_xx_010_110_xxx_1_x_xx;
      patterns[8459] = 33'b0100111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8460] = 33'b0000011000111110_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8461] = 33'b0000111000111110_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8462] = 33'b0000111000111110_0_0_00_000_000_000_0_0_00;
      patterns[8463] = 33'b1000011000100011_0_1_00_010_011_110_0_x_00;
      patterns[8464] = 33'b1000111000100011_1_1_00_010_011_110_0_x_00;
      patterns[8465] = 33'b1000111000100011_0_0_00_000_000_000_0_0_00;
      patterns[8466] = 33'b1001011000100011_0_1_01_010_011_110_0_x_00;
      patterns[8467] = 33'b1001111000100011_1_1_01_010_011_110_0_x_00;
      patterns[8468] = 33'b1001111000100011_0_0_00_000_000_000_0_0_00;
      patterns[8469] = 33'b1010011000100011_0_1_10_010_011_110_0_x_00;
      patterns[8470] = 33'b1010111000100011_1_1_10_010_011_110_0_x_00;
      patterns[8471] = 33'b1010111000100011_0_0_00_000_000_000_0_0_00;
      patterns[8472] = 33'b1011011000100011_0_1_11_010_011_110_0_x_00;
      patterns[8473] = 33'b1011111000100011_1_1_11_010_011_110_0_x_00;
      patterns[8474] = 33'b1011111000100011_0_0_00_000_000_000_0_0_00;
      patterns[8475] = 33'b0101011000100000_0_1_xx_010_xxx_110_0_1_01;
      patterns[8476] = 33'b0101111000100000_1_1_xx_010_xxx_110_0_1_01;
      patterns[8477] = 33'b0101111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8478] = 33'b0100011000100000_0_0_xx_010_110_xxx_1_x_xx;
      patterns[8479] = 33'b0100111000100000_1_0_xx_010_110_xxx_1_x_xx;
      patterns[8480] = 33'b0100111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8481] = 33'b0000011010101011_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8482] = 33'b0000111010101011_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8483] = 33'b0000111010101011_0_0_00_000_000_000_0_0_00;
      patterns[8484] = 33'b1000011000100100_0_1_00_010_100_110_0_x_00;
      patterns[8485] = 33'b1000111000100100_1_1_00_010_100_110_0_x_00;
      patterns[8486] = 33'b1000111000100100_0_0_00_000_000_000_0_0_00;
      patterns[8487] = 33'b1001011000100100_0_1_01_010_100_110_0_x_00;
      patterns[8488] = 33'b1001111000100100_1_1_01_010_100_110_0_x_00;
      patterns[8489] = 33'b1001111000100100_0_0_00_000_000_000_0_0_00;
      patterns[8490] = 33'b1010011000100100_0_1_10_010_100_110_0_x_00;
      patterns[8491] = 33'b1010111000100100_1_1_10_010_100_110_0_x_00;
      patterns[8492] = 33'b1010111000100100_0_0_00_000_000_000_0_0_00;
      patterns[8493] = 33'b1011011000100100_0_1_11_010_100_110_0_x_00;
      patterns[8494] = 33'b1011111000100100_1_1_11_010_100_110_0_x_00;
      patterns[8495] = 33'b1011111000100100_0_0_00_000_000_000_0_0_00;
      patterns[8496] = 33'b0101011000100000_0_1_xx_010_xxx_110_0_1_01;
      patterns[8497] = 33'b0101111000100000_1_1_xx_010_xxx_110_0_1_01;
      patterns[8498] = 33'b0101111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8499] = 33'b0100011000100000_0_0_xx_010_110_xxx_1_x_xx;
      patterns[8500] = 33'b0100111000100000_1_0_xx_010_110_xxx_1_x_xx;
      patterns[8501] = 33'b0100111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8502] = 33'b0000011010011001_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8503] = 33'b0000111010011001_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8504] = 33'b0000111010011001_0_0_00_000_000_000_0_0_00;
      patterns[8505] = 33'b1000011000100101_0_1_00_010_101_110_0_x_00;
      patterns[8506] = 33'b1000111000100101_1_1_00_010_101_110_0_x_00;
      patterns[8507] = 33'b1000111000100101_0_0_00_000_000_000_0_0_00;
      patterns[8508] = 33'b1001011000100101_0_1_01_010_101_110_0_x_00;
      patterns[8509] = 33'b1001111000100101_1_1_01_010_101_110_0_x_00;
      patterns[8510] = 33'b1001111000100101_0_0_00_000_000_000_0_0_00;
      patterns[8511] = 33'b1010011000100101_0_1_10_010_101_110_0_x_00;
      patterns[8512] = 33'b1010111000100101_1_1_10_010_101_110_0_x_00;
      patterns[8513] = 33'b1010111000100101_0_0_00_000_000_000_0_0_00;
      patterns[8514] = 33'b1011011000100101_0_1_11_010_101_110_0_x_00;
      patterns[8515] = 33'b1011111000100101_1_1_11_010_101_110_0_x_00;
      patterns[8516] = 33'b1011111000100101_0_0_00_000_000_000_0_0_00;
      patterns[8517] = 33'b0101011000100000_0_1_xx_010_xxx_110_0_1_01;
      patterns[8518] = 33'b0101111000100000_1_1_xx_010_xxx_110_0_1_01;
      patterns[8519] = 33'b0101111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8520] = 33'b0100011000100000_0_0_xx_010_110_xxx_1_x_xx;
      patterns[8521] = 33'b0100111000100000_1_0_xx_010_110_xxx_1_x_xx;
      patterns[8522] = 33'b0100111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8523] = 33'b0000011001101001_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8524] = 33'b0000111001101001_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8525] = 33'b0000111001101001_0_0_00_000_000_000_0_0_00;
      patterns[8526] = 33'b1000011000100110_0_1_00_010_110_110_0_x_00;
      patterns[8527] = 33'b1000111000100110_1_1_00_010_110_110_0_x_00;
      patterns[8528] = 33'b1000111000100110_0_0_00_000_000_000_0_0_00;
      patterns[8529] = 33'b1001011000100110_0_1_01_010_110_110_0_x_00;
      patterns[8530] = 33'b1001111000100110_1_1_01_010_110_110_0_x_00;
      patterns[8531] = 33'b1001111000100110_0_0_00_000_000_000_0_0_00;
      patterns[8532] = 33'b1010011000100110_0_1_10_010_110_110_0_x_00;
      patterns[8533] = 33'b1010111000100110_1_1_10_010_110_110_0_x_00;
      patterns[8534] = 33'b1010111000100110_0_0_00_000_000_000_0_0_00;
      patterns[8535] = 33'b1011011000100110_0_1_11_010_110_110_0_x_00;
      patterns[8536] = 33'b1011111000100110_1_1_11_010_110_110_0_x_00;
      patterns[8537] = 33'b1011111000100110_0_0_00_000_000_000_0_0_00;
      patterns[8538] = 33'b0101011000100000_0_1_xx_010_xxx_110_0_1_01;
      patterns[8539] = 33'b0101111000100000_1_1_xx_010_xxx_110_0_1_01;
      patterns[8540] = 33'b0101111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8541] = 33'b0100011000100000_0_0_xx_010_110_xxx_1_x_xx;
      patterns[8542] = 33'b0100111000100000_1_0_xx_010_110_xxx_1_x_xx;
      patterns[8543] = 33'b0100111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8544] = 33'b0000011001101100_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8545] = 33'b0000111001101100_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8546] = 33'b0000111001101100_0_0_00_000_000_000_0_0_00;
      patterns[8547] = 33'b1000011000100111_0_1_00_010_111_110_0_x_00;
      patterns[8548] = 33'b1000111000100111_1_1_00_010_111_110_0_x_00;
      patterns[8549] = 33'b1000111000100111_0_0_00_000_000_000_0_0_00;
      patterns[8550] = 33'b1001011000100111_0_1_01_010_111_110_0_x_00;
      patterns[8551] = 33'b1001111000100111_1_1_01_010_111_110_0_x_00;
      patterns[8552] = 33'b1001111000100111_0_0_00_000_000_000_0_0_00;
      patterns[8553] = 33'b1010011000100111_0_1_10_010_111_110_0_x_00;
      patterns[8554] = 33'b1010111000100111_1_1_10_010_111_110_0_x_00;
      patterns[8555] = 33'b1010111000100111_0_0_00_000_000_000_0_0_00;
      patterns[8556] = 33'b1011011000100111_0_1_11_010_111_110_0_x_00;
      patterns[8557] = 33'b1011111000100111_1_1_11_010_111_110_0_x_00;
      patterns[8558] = 33'b1011111000100111_0_0_00_000_000_000_0_0_00;
      patterns[8559] = 33'b0101011000100000_0_1_xx_010_xxx_110_0_1_01;
      patterns[8560] = 33'b0101111000100000_1_1_xx_010_xxx_110_0_1_01;
      patterns[8561] = 33'b0101111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8562] = 33'b0100011000100000_0_0_xx_010_110_xxx_1_x_xx;
      patterns[8563] = 33'b0100111000100000_1_0_xx_010_110_xxx_1_x_xx;
      patterns[8564] = 33'b0100111000100000_0_0_00_000_000_000_0_0_00;
      patterns[8565] = 33'b0000011011010110_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8566] = 33'b0000111011010110_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8567] = 33'b0000111011010110_0_0_00_000_000_000_0_0_00;
      patterns[8568] = 33'b1000011000110000_0_1_00_011_000_110_0_x_00;
      patterns[8569] = 33'b1000111000110000_1_1_00_011_000_110_0_x_00;
      patterns[8570] = 33'b1000111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8571] = 33'b1001011000110000_0_1_01_011_000_110_0_x_00;
      patterns[8572] = 33'b1001111000110000_1_1_01_011_000_110_0_x_00;
      patterns[8573] = 33'b1001111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8574] = 33'b1010011000110000_0_1_10_011_000_110_0_x_00;
      patterns[8575] = 33'b1010111000110000_1_1_10_011_000_110_0_x_00;
      patterns[8576] = 33'b1010111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8577] = 33'b1011011000110000_0_1_11_011_000_110_0_x_00;
      patterns[8578] = 33'b1011111000110000_1_1_11_011_000_110_0_x_00;
      patterns[8579] = 33'b1011111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8580] = 33'b0101011000110000_0_1_xx_011_xxx_110_0_1_01;
      patterns[8581] = 33'b0101111000110000_1_1_xx_011_xxx_110_0_1_01;
      patterns[8582] = 33'b0101111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8583] = 33'b0100011000110000_0_0_xx_011_110_xxx_1_x_xx;
      patterns[8584] = 33'b0100111000110000_1_0_xx_011_110_xxx_1_x_xx;
      patterns[8585] = 33'b0100111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8586] = 33'b0000011010010111_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8587] = 33'b0000111010010111_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8588] = 33'b0000111010010111_0_0_00_000_000_000_0_0_00;
      patterns[8589] = 33'b1000011000110001_0_1_00_011_001_110_0_x_00;
      patterns[8590] = 33'b1000111000110001_1_1_00_011_001_110_0_x_00;
      patterns[8591] = 33'b1000111000110001_0_0_00_000_000_000_0_0_00;
      patterns[8592] = 33'b1001011000110001_0_1_01_011_001_110_0_x_00;
      patterns[8593] = 33'b1001111000110001_1_1_01_011_001_110_0_x_00;
      patterns[8594] = 33'b1001111000110001_0_0_00_000_000_000_0_0_00;
      patterns[8595] = 33'b1010011000110001_0_1_10_011_001_110_0_x_00;
      patterns[8596] = 33'b1010111000110001_1_1_10_011_001_110_0_x_00;
      patterns[8597] = 33'b1010111000110001_0_0_00_000_000_000_0_0_00;
      patterns[8598] = 33'b1011011000110001_0_1_11_011_001_110_0_x_00;
      patterns[8599] = 33'b1011111000110001_1_1_11_011_001_110_0_x_00;
      patterns[8600] = 33'b1011111000110001_0_0_00_000_000_000_0_0_00;
      patterns[8601] = 33'b0101011000110000_0_1_xx_011_xxx_110_0_1_01;
      patterns[8602] = 33'b0101111000110000_1_1_xx_011_xxx_110_0_1_01;
      patterns[8603] = 33'b0101111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8604] = 33'b0100011000110000_0_0_xx_011_110_xxx_1_x_xx;
      patterns[8605] = 33'b0100111000110000_1_0_xx_011_110_xxx_1_x_xx;
      patterns[8606] = 33'b0100111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8607] = 33'b0000011001110110_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8608] = 33'b0000111001110110_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8609] = 33'b0000111001110110_0_0_00_000_000_000_0_0_00;
      patterns[8610] = 33'b1000011000110010_0_1_00_011_010_110_0_x_00;
      patterns[8611] = 33'b1000111000110010_1_1_00_011_010_110_0_x_00;
      patterns[8612] = 33'b1000111000110010_0_0_00_000_000_000_0_0_00;
      patterns[8613] = 33'b1001011000110010_0_1_01_011_010_110_0_x_00;
      patterns[8614] = 33'b1001111000110010_1_1_01_011_010_110_0_x_00;
      patterns[8615] = 33'b1001111000110010_0_0_00_000_000_000_0_0_00;
      patterns[8616] = 33'b1010011000110010_0_1_10_011_010_110_0_x_00;
      patterns[8617] = 33'b1010111000110010_1_1_10_011_010_110_0_x_00;
      patterns[8618] = 33'b1010111000110010_0_0_00_000_000_000_0_0_00;
      patterns[8619] = 33'b1011011000110010_0_1_11_011_010_110_0_x_00;
      patterns[8620] = 33'b1011111000110010_1_1_11_011_010_110_0_x_00;
      patterns[8621] = 33'b1011111000110010_0_0_00_000_000_000_0_0_00;
      patterns[8622] = 33'b0101011000110000_0_1_xx_011_xxx_110_0_1_01;
      patterns[8623] = 33'b0101111000110000_1_1_xx_011_xxx_110_0_1_01;
      patterns[8624] = 33'b0101111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8625] = 33'b0100011000110000_0_0_xx_011_110_xxx_1_x_xx;
      patterns[8626] = 33'b0100111000110000_1_0_xx_011_110_xxx_1_x_xx;
      patterns[8627] = 33'b0100111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8628] = 33'b0000011001111011_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8629] = 33'b0000111001111011_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8630] = 33'b0000111001111011_0_0_00_000_000_000_0_0_00;
      patterns[8631] = 33'b1000011000110011_0_1_00_011_011_110_0_x_00;
      patterns[8632] = 33'b1000111000110011_1_1_00_011_011_110_0_x_00;
      patterns[8633] = 33'b1000111000110011_0_0_00_000_000_000_0_0_00;
      patterns[8634] = 33'b1001011000110011_0_1_01_011_011_110_0_x_00;
      patterns[8635] = 33'b1001111000110011_1_1_01_011_011_110_0_x_00;
      patterns[8636] = 33'b1001111000110011_0_0_00_000_000_000_0_0_00;
      patterns[8637] = 33'b1010011000110011_0_1_10_011_011_110_0_x_00;
      patterns[8638] = 33'b1010111000110011_1_1_10_011_011_110_0_x_00;
      patterns[8639] = 33'b1010111000110011_0_0_00_000_000_000_0_0_00;
      patterns[8640] = 33'b1011011000110011_0_1_11_011_011_110_0_x_00;
      patterns[8641] = 33'b1011111000110011_1_1_11_011_011_110_0_x_00;
      patterns[8642] = 33'b1011111000110011_0_0_00_000_000_000_0_0_00;
      patterns[8643] = 33'b0101011000110000_0_1_xx_011_xxx_110_0_1_01;
      patterns[8644] = 33'b0101111000110000_1_1_xx_011_xxx_110_0_1_01;
      patterns[8645] = 33'b0101111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8646] = 33'b0100011000110000_0_0_xx_011_110_xxx_1_x_xx;
      patterns[8647] = 33'b0100111000110000_1_0_xx_011_110_xxx_1_x_xx;
      patterns[8648] = 33'b0100111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8649] = 33'b0000011000111111_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8650] = 33'b0000111000111111_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8651] = 33'b0000111000111111_0_0_00_000_000_000_0_0_00;
      patterns[8652] = 33'b1000011000110100_0_1_00_011_100_110_0_x_00;
      patterns[8653] = 33'b1000111000110100_1_1_00_011_100_110_0_x_00;
      patterns[8654] = 33'b1000111000110100_0_0_00_000_000_000_0_0_00;
      patterns[8655] = 33'b1001011000110100_0_1_01_011_100_110_0_x_00;
      patterns[8656] = 33'b1001111000110100_1_1_01_011_100_110_0_x_00;
      patterns[8657] = 33'b1001111000110100_0_0_00_000_000_000_0_0_00;
      patterns[8658] = 33'b1010011000110100_0_1_10_011_100_110_0_x_00;
      patterns[8659] = 33'b1010111000110100_1_1_10_011_100_110_0_x_00;
      patterns[8660] = 33'b1010111000110100_0_0_00_000_000_000_0_0_00;
      patterns[8661] = 33'b1011011000110100_0_1_11_011_100_110_0_x_00;
      patterns[8662] = 33'b1011111000110100_1_1_11_011_100_110_0_x_00;
      patterns[8663] = 33'b1011111000110100_0_0_00_000_000_000_0_0_00;
      patterns[8664] = 33'b0101011000110000_0_1_xx_011_xxx_110_0_1_01;
      patterns[8665] = 33'b0101111000110000_1_1_xx_011_xxx_110_0_1_01;
      patterns[8666] = 33'b0101111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8667] = 33'b0100011000110000_0_0_xx_011_110_xxx_1_x_xx;
      patterns[8668] = 33'b0100111000110000_1_0_xx_011_110_xxx_1_x_xx;
      patterns[8669] = 33'b0100111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8670] = 33'b0000011001101011_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8671] = 33'b0000111001101011_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8672] = 33'b0000111001101011_0_0_00_000_000_000_0_0_00;
      patterns[8673] = 33'b1000011000110101_0_1_00_011_101_110_0_x_00;
      patterns[8674] = 33'b1000111000110101_1_1_00_011_101_110_0_x_00;
      patterns[8675] = 33'b1000111000110101_0_0_00_000_000_000_0_0_00;
      patterns[8676] = 33'b1001011000110101_0_1_01_011_101_110_0_x_00;
      patterns[8677] = 33'b1001111000110101_1_1_01_011_101_110_0_x_00;
      patterns[8678] = 33'b1001111000110101_0_0_00_000_000_000_0_0_00;
      patterns[8679] = 33'b1010011000110101_0_1_10_011_101_110_0_x_00;
      patterns[8680] = 33'b1010111000110101_1_1_10_011_101_110_0_x_00;
      patterns[8681] = 33'b1010111000110101_0_0_00_000_000_000_0_0_00;
      patterns[8682] = 33'b1011011000110101_0_1_11_011_101_110_0_x_00;
      patterns[8683] = 33'b1011111000110101_1_1_11_011_101_110_0_x_00;
      patterns[8684] = 33'b1011111000110101_0_0_00_000_000_000_0_0_00;
      patterns[8685] = 33'b0101011000110000_0_1_xx_011_xxx_110_0_1_01;
      patterns[8686] = 33'b0101111000110000_1_1_xx_011_xxx_110_0_1_01;
      patterns[8687] = 33'b0101111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8688] = 33'b0100011000110000_0_0_xx_011_110_xxx_1_x_xx;
      patterns[8689] = 33'b0100111000110000_1_0_xx_011_110_xxx_1_x_xx;
      patterns[8690] = 33'b0100111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8691] = 33'b0000011000111100_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8692] = 33'b0000111000111100_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8693] = 33'b0000111000111100_0_0_00_000_000_000_0_0_00;
      patterns[8694] = 33'b1000011000110110_0_1_00_011_110_110_0_x_00;
      patterns[8695] = 33'b1000111000110110_1_1_00_011_110_110_0_x_00;
      patterns[8696] = 33'b1000111000110110_0_0_00_000_000_000_0_0_00;
      patterns[8697] = 33'b1001011000110110_0_1_01_011_110_110_0_x_00;
      patterns[8698] = 33'b1001111000110110_1_1_01_011_110_110_0_x_00;
      patterns[8699] = 33'b1001111000110110_0_0_00_000_000_000_0_0_00;
      patterns[8700] = 33'b1010011000110110_0_1_10_011_110_110_0_x_00;
      patterns[8701] = 33'b1010111000110110_1_1_10_011_110_110_0_x_00;
      patterns[8702] = 33'b1010111000110110_0_0_00_000_000_000_0_0_00;
      patterns[8703] = 33'b1011011000110110_0_1_11_011_110_110_0_x_00;
      patterns[8704] = 33'b1011111000110110_1_1_11_011_110_110_0_x_00;
      patterns[8705] = 33'b1011111000110110_0_0_00_000_000_000_0_0_00;
      patterns[8706] = 33'b0101011000110000_0_1_xx_011_xxx_110_0_1_01;
      patterns[8707] = 33'b0101111000110000_1_1_xx_011_xxx_110_0_1_01;
      patterns[8708] = 33'b0101111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8709] = 33'b0100011000110000_0_0_xx_011_110_xxx_1_x_xx;
      patterns[8710] = 33'b0100111000110000_1_0_xx_011_110_xxx_1_x_xx;
      patterns[8711] = 33'b0100111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8712] = 33'b0000011010100100_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8713] = 33'b0000111010100100_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8714] = 33'b0000111010100100_0_0_00_000_000_000_0_0_00;
      patterns[8715] = 33'b1000011000110111_0_1_00_011_111_110_0_x_00;
      patterns[8716] = 33'b1000111000110111_1_1_00_011_111_110_0_x_00;
      patterns[8717] = 33'b1000111000110111_0_0_00_000_000_000_0_0_00;
      patterns[8718] = 33'b1001011000110111_0_1_01_011_111_110_0_x_00;
      patterns[8719] = 33'b1001111000110111_1_1_01_011_111_110_0_x_00;
      patterns[8720] = 33'b1001111000110111_0_0_00_000_000_000_0_0_00;
      patterns[8721] = 33'b1010011000110111_0_1_10_011_111_110_0_x_00;
      patterns[8722] = 33'b1010111000110111_1_1_10_011_111_110_0_x_00;
      patterns[8723] = 33'b1010111000110111_0_0_00_000_000_000_0_0_00;
      patterns[8724] = 33'b1011011000110111_0_1_11_011_111_110_0_x_00;
      patterns[8725] = 33'b1011111000110111_1_1_11_011_111_110_0_x_00;
      patterns[8726] = 33'b1011111000110111_0_0_00_000_000_000_0_0_00;
      patterns[8727] = 33'b0101011000110000_0_1_xx_011_xxx_110_0_1_01;
      patterns[8728] = 33'b0101111000110000_1_1_xx_011_xxx_110_0_1_01;
      patterns[8729] = 33'b0101111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8730] = 33'b0100011000110000_0_0_xx_011_110_xxx_1_x_xx;
      patterns[8731] = 33'b0100111000110000_1_0_xx_011_110_xxx_1_x_xx;
      patterns[8732] = 33'b0100111000110000_0_0_00_000_000_000_0_0_00;
      patterns[8733] = 33'b0000011001010110_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8734] = 33'b0000111001010110_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8735] = 33'b0000111001010110_0_0_00_000_000_000_0_0_00;
      patterns[8736] = 33'b1000011001000000_0_1_00_100_000_110_0_x_00;
      patterns[8737] = 33'b1000111001000000_1_1_00_100_000_110_0_x_00;
      patterns[8738] = 33'b1000111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8739] = 33'b1001011001000000_0_1_01_100_000_110_0_x_00;
      patterns[8740] = 33'b1001111001000000_1_1_01_100_000_110_0_x_00;
      patterns[8741] = 33'b1001111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8742] = 33'b1010011001000000_0_1_10_100_000_110_0_x_00;
      patterns[8743] = 33'b1010111001000000_1_1_10_100_000_110_0_x_00;
      patterns[8744] = 33'b1010111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8745] = 33'b1011011001000000_0_1_11_100_000_110_0_x_00;
      patterns[8746] = 33'b1011111001000000_1_1_11_100_000_110_0_x_00;
      patterns[8747] = 33'b1011111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8748] = 33'b0101011001000000_0_1_xx_100_xxx_110_0_1_01;
      patterns[8749] = 33'b0101111001000000_1_1_xx_100_xxx_110_0_1_01;
      patterns[8750] = 33'b0101111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8751] = 33'b0100011001000000_0_0_xx_100_110_xxx_1_x_xx;
      patterns[8752] = 33'b0100111001000000_1_0_xx_100_110_xxx_1_x_xx;
      patterns[8753] = 33'b0100111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8754] = 33'b0000011010110000_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8755] = 33'b0000111010110000_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8756] = 33'b0000111010110000_0_0_00_000_000_000_0_0_00;
      patterns[8757] = 33'b1000011001000001_0_1_00_100_001_110_0_x_00;
      patterns[8758] = 33'b1000111001000001_1_1_00_100_001_110_0_x_00;
      patterns[8759] = 33'b1000111001000001_0_0_00_000_000_000_0_0_00;
      patterns[8760] = 33'b1001011001000001_0_1_01_100_001_110_0_x_00;
      patterns[8761] = 33'b1001111001000001_1_1_01_100_001_110_0_x_00;
      patterns[8762] = 33'b1001111001000001_0_0_00_000_000_000_0_0_00;
      patterns[8763] = 33'b1010011001000001_0_1_10_100_001_110_0_x_00;
      patterns[8764] = 33'b1010111001000001_1_1_10_100_001_110_0_x_00;
      patterns[8765] = 33'b1010111001000001_0_0_00_000_000_000_0_0_00;
      patterns[8766] = 33'b1011011001000001_0_1_11_100_001_110_0_x_00;
      patterns[8767] = 33'b1011111001000001_1_1_11_100_001_110_0_x_00;
      patterns[8768] = 33'b1011111001000001_0_0_00_000_000_000_0_0_00;
      patterns[8769] = 33'b0101011001000000_0_1_xx_100_xxx_110_0_1_01;
      patterns[8770] = 33'b0101111001000000_1_1_xx_100_xxx_110_0_1_01;
      patterns[8771] = 33'b0101111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8772] = 33'b0100011001000000_0_0_xx_100_110_xxx_1_x_xx;
      patterns[8773] = 33'b0100111001000000_1_0_xx_100_110_xxx_1_x_xx;
      patterns[8774] = 33'b0100111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8775] = 33'b0000011011101010_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8776] = 33'b0000111011101010_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8777] = 33'b0000111011101010_0_0_00_000_000_000_0_0_00;
      patterns[8778] = 33'b1000011001000010_0_1_00_100_010_110_0_x_00;
      patterns[8779] = 33'b1000111001000010_1_1_00_100_010_110_0_x_00;
      patterns[8780] = 33'b1000111001000010_0_0_00_000_000_000_0_0_00;
      patterns[8781] = 33'b1001011001000010_0_1_01_100_010_110_0_x_00;
      patterns[8782] = 33'b1001111001000010_1_1_01_100_010_110_0_x_00;
      patterns[8783] = 33'b1001111001000010_0_0_00_000_000_000_0_0_00;
      patterns[8784] = 33'b1010011001000010_0_1_10_100_010_110_0_x_00;
      patterns[8785] = 33'b1010111001000010_1_1_10_100_010_110_0_x_00;
      patterns[8786] = 33'b1010111001000010_0_0_00_000_000_000_0_0_00;
      patterns[8787] = 33'b1011011001000010_0_1_11_100_010_110_0_x_00;
      patterns[8788] = 33'b1011111001000010_1_1_11_100_010_110_0_x_00;
      patterns[8789] = 33'b1011111001000010_0_0_00_000_000_000_0_0_00;
      patterns[8790] = 33'b0101011001000000_0_1_xx_100_xxx_110_0_1_01;
      patterns[8791] = 33'b0101111001000000_1_1_xx_100_xxx_110_0_1_01;
      patterns[8792] = 33'b0101111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8793] = 33'b0100011001000000_0_0_xx_100_110_xxx_1_x_xx;
      patterns[8794] = 33'b0100111001000000_1_0_xx_100_110_xxx_1_x_xx;
      patterns[8795] = 33'b0100111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8796] = 33'b0000011010100000_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8797] = 33'b0000111010100000_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8798] = 33'b0000111010100000_0_0_00_000_000_000_0_0_00;
      patterns[8799] = 33'b1000011001000011_0_1_00_100_011_110_0_x_00;
      patterns[8800] = 33'b1000111001000011_1_1_00_100_011_110_0_x_00;
      patterns[8801] = 33'b1000111001000011_0_0_00_000_000_000_0_0_00;
      patterns[8802] = 33'b1001011001000011_0_1_01_100_011_110_0_x_00;
      patterns[8803] = 33'b1001111001000011_1_1_01_100_011_110_0_x_00;
      patterns[8804] = 33'b1001111001000011_0_0_00_000_000_000_0_0_00;
      patterns[8805] = 33'b1010011001000011_0_1_10_100_011_110_0_x_00;
      patterns[8806] = 33'b1010111001000011_1_1_10_100_011_110_0_x_00;
      patterns[8807] = 33'b1010111001000011_0_0_00_000_000_000_0_0_00;
      patterns[8808] = 33'b1011011001000011_0_1_11_100_011_110_0_x_00;
      patterns[8809] = 33'b1011111001000011_1_1_11_100_011_110_0_x_00;
      patterns[8810] = 33'b1011111001000011_0_0_00_000_000_000_0_0_00;
      patterns[8811] = 33'b0101011001000000_0_1_xx_100_xxx_110_0_1_01;
      patterns[8812] = 33'b0101111001000000_1_1_xx_100_xxx_110_0_1_01;
      patterns[8813] = 33'b0101111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8814] = 33'b0100011001000000_0_0_xx_100_110_xxx_1_x_xx;
      patterns[8815] = 33'b0100111001000000_1_0_xx_100_110_xxx_1_x_xx;
      patterns[8816] = 33'b0100111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8817] = 33'b0000011011010010_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8818] = 33'b0000111011010010_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8819] = 33'b0000111011010010_0_0_00_000_000_000_0_0_00;
      patterns[8820] = 33'b1000011001000100_0_1_00_100_100_110_0_x_00;
      patterns[8821] = 33'b1000111001000100_1_1_00_100_100_110_0_x_00;
      patterns[8822] = 33'b1000111001000100_0_0_00_000_000_000_0_0_00;
      patterns[8823] = 33'b1001011001000100_0_1_01_100_100_110_0_x_00;
      patterns[8824] = 33'b1001111001000100_1_1_01_100_100_110_0_x_00;
      patterns[8825] = 33'b1001111001000100_0_0_00_000_000_000_0_0_00;
      patterns[8826] = 33'b1010011001000100_0_1_10_100_100_110_0_x_00;
      patterns[8827] = 33'b1010111001000100_1_1_10_100_100_110_0_x_00;
      patterns[8828] = 33'b1010111001000100_0_0_00_000_000_000_0_0_00;
      patterns[8829] = 33'b1011011001000100_0_1_11_100_100_110_0_x_00;
      patterns[8830] = 33'b1011111001000100_1_1_11_100_100_110_0_x_00;
      patterns[8831] = 33'b1011111001000100_0_0_00_000_000_000_0_0_00;
      patterns[8832] = 33'b0101011001000000_0_1_xx_100_xxx_110_0_1_01;
      patterns[8833] = 33'b0101111001000000_1_1_xx_100_xxx_110_0_1_01;
      patterns[8834] = 33'b0101111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8835] = 33'b0100011001000000_0_0_xx_100_110_xxx_1_x_xx;
      patterns[8836] = 33'b0100111001000000_1_0_xx_100_110_xxx_1_x_xx;
      patterns[8837] = 33'b0100111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8838] = 33'b0000011001111000_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8839] = 33'b0000111001111000_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8840] = 33'b0000111001111000_0_0_00_000_000_000_0_0_00;
      patterns[8841] = 33'b1000011001000101_0_1_00_100_101_110_0_x_00;
      patterns[8842] = 33'b1000111001000101_1_1_00_100_101_110_0_x_00;
      patterns[8843] = 33'b1000111001000101_0_0_00_000_000_000_0_0_00;
      patterns[8844] = 33'b1001011001000101_0_1_01_100_101_110_0_x_00;
      patterns[8845] = 33'b1001111001000101_1_1_01_100_101_110_0_x_00;
      patterns[8846] = 33'b1001111001000101_0_0_00_000_000_000_0_0_00;
      patterns[8847] = 33'b1010011001000101_0_1_10_100_101_110_0_x_00;
      patterns[8848] = 33'b1010111001000101_1_1_10_100_101_110_0_x_00;
      patterns[8849] = 33'b1010111001000101_0_0_00_000_000_000_0_0_00;
      patterns[8850] = 33'b1011011001000101_0_1_11_100_101_110_0_x_00;
      patterns[8851] = 33'b1011111001000101_1_1_11_100_101_110_0_x_00;
      patterns[8852] = 33'b1011111001000101_0_0_00_000_000_000_0_0_00;
      patterns[8853] = 33'b0101011001000000_0_1_xx_100_xxx_110_0_1_01;
      patterns[8854] = 33'b0101111001000000_1_1_xx_100_xxx_110_0_1_01;
      patterns[8855] = 33'b0101111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8856] = 33'b0100011001000000_0_0_xx_100_110_xxx_1_x_xx;
      patterns[8857] = 33'b0100111001000000_1_0_xx_100_110_xxx_1_x_xx;
      patterns[8858] = 33'b0100111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8859] = 33'b0000011000010000_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8860] = 33'b0000111000010000_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8861] = 33'b0000111000010000_0_0_00_000_000_000_0_0_00;
      patterns[8862] = 33'b1000011001000110_0_1_00_100_110_110_0_x_00;
      patterns[8863] = 33'b1000111001000110_1_1_00_100_110_110_0_x_00;
      patterns[8864] = 33'b1000111001000110_0_0_00_000_000_000_0_0_00;
      patterns[8865] = 33'b1001011001000110_0_1_01_100_110_110_0_x_00;
      patterns[8866] = 33'b1001111001000110_1_1_01_100_110_110_0_x_00;
      patterns[8867] = 33'b1001111001000110_0_0_00_000_000_000_0_0_00;
      patterns[8868] = 33'b1010011001000110_0_1_10_100_110_110_0_x_00;
      patterns[8869] = 33'b1010111001000110_1_1_10_100_110_110_0_x_00;
      patterns[8870] = 33'b1010111001000110_0_0_00_000_000_000_0_0_00;
      patterns[8871] = 33'b1011011001000110_0_1_11_100_110_110_0_x_00;
      patterns[8872] = 33'b1011111001000110_1_1_11_100_110_110_0_x_00;
      patterns[8873] = 33'b1011111001000110_0_0_00_000_000_000_0_0_00;
      patterns[8874] = 33'b0101011001000000_0_1_xx_100_xxx_110_0_1_01;
      patterns[8875] = 33'b0101111001000000_1_1_xx_100_xxx_110_0_1_01;
      patterns[8876] = 33'b0101111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8877] = 33'b0100011001000000_0_0_xx_100_110_xxx_1_x_xx;
      patterns[8878] = 33'b0100111001000000_1_0_xx_100_110_xxx_1_x_xx;
      patterns[8879] = 33'b0100111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8880] = 33'b0000011001011000_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8881] = 33'b0000111001011000_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8882] = 33'b0000111001011000_0_0_00_000_000_000_0_0_00;
      patterns[8883] = 33'b1000011001000111_0_1_00_100_111_110_0_x_00;
      patterns[8884] = 33'b1000111001000111_1_1_00_100_111_110_0_x_00;
      patterns[8885] = 33'b1000111001000111_0_0_00_000_000_000_0_0_00;
      patterns[8886] = 33'b1001011001000111_0_1_01_100_111_110_0_x_00;
      patterns[8887] = 33'b1001111001000111_1_1_01_100_111_110_0_x_00;
      patterns[8888] = 33'b1001111001000111_0_0_00_000_000_000_0_0_00;
      patterns[8889] = 33'b1010011001000111_0_1_10_100_111_110_0_x_00;
      patterns[8890] = 33'b1010111001000111_1_1_10_100_111_110_0_x_00;
      patterns[8891] = 33'b1010111001000111_0_0_00_000_000_000_0_0_00;
      patterns[8892] = 33'b1011011001000111_0_1_11_100_111_110_0_x_00;
      patterns[8893] = 33'b1011111001000111_1_1_11_100_111_110_0_x_00;
      patterns[8894] = 33'b1011111001000111_0_0_00_000_000_000_0_0_00;
      patterns[8895] = 33'b0101011001000000_0_1_xx_100_xxx_110_0_1_01;
      patterns[8896] = 33'b0101111001000000_1_1_xx_100_xxx_110_0_1_01;
      patterns[8897] = 33'b0101111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8898] = 33'b0100011001000000_0_0_xx_100_110_xxx_1_x_xx;
      patterns[8899] = 33'b0100111001000000_1_0_xx_100_110_xxx_1_x_xx;
      patterns[8900] = 33'b0100111001000000_0_0_00_000_000_000_0_0_00;
      patterns[8901] = 33'b0000011011111001_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8902] = 33'b0000111011111001_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8903] = 33'b0000111011111001_0_0_00_000_000_000_0_0_00;
      patterns[8904] = 33'b1000011001010000_0_1_00_101_000_110_0_x_00;
      patterns[8905] = 33'b1000111001010000_1_1_00_101_000_110_0_x_00;
      patterns[8906] = 33'b1000111001010000_0_0_00_000_000_000_0_0_00;
      patterns[8907] = 33'b1001011001010000_0_1_01_101_000_110_0_x_00;
      patterns[8908] = 33'b1001111001010000_1_1_01_101_000_110_0_x_00;
      patterns[8909] = 33'b1001111001010000_0_0_00_000_000_000_0_0_00;
      patterns[8910] = 33'b1010011001010000_0_1_10_101_000_110_0_x_00;
      patterns[8911] = 33'b1010111001010000_1_1_10_101_000_110_0_x_00;
      patterns[8912] = 33'b1010111001010000_0_0_00_000_000_000_0_0_00;
      patterns[8913] = 33'b1011011001010000_0_1_11_101_000_110_0_x_00;
      patterns[8914] = 33'b1011111001010000_1_1_11_101_000_110_0_x_00;
      patterns[8915] = 33'b1011111001010000_0_0_00_000_000_000_0_0_00;
      patterns[8916] = 33'b0101011001010000_0_1_xx_101_xxx_110_0_1_01;
      patterns[8917] = 33'b0101111001010000_1_1_xx_101_xxx_110_0_1_01;
      patterns[8918] = 33'b0101111001010000_0_0_00_000_000_000_0_0_00;
      patterns[8919] = 33'b0100011001010000_0_0_xx_101_110_xxx_1_x_xx;
      patterns[8920] = 33'b0100111001010000_1_0_xx_101_110_xxx_1_x_xx;
      patterns[8921] = 33'b0100111001010000_0_0_00_000_000_000_0_0_00;
      patterns[8922] = 33'b0000011000011010_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8923] = 33'b0000111000011010_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8924] = 33'b0000111000011010_0_0_00_000_000_000_0_0_00;
      patterns[8925] = 33'b1000011001010001_0_1_00_101_001_110_0_x_00;
      patterns[8926] = 33'b1000111001010001_1_1_00_101_001_110_0_x_00;
      patterns[8927] = 33'b1000111001010001_0_0_00_000_000_000_0_0_00;
      patterns[8928] = 33'b1001011001010001_0_1_01_101_001_110_0_x_00;
      patterns[8929] = 33'b1001111001010001_1_1_01_101_001_110_0_x_00;
      patterns[8930] = 33'b1001111001010001_0_0_00_000_000_000_0_0_00;
      patterns[8931] = 33'b1010011001010001_0_1_10_101_001_110_0_x_00;
      patterns[8932] = 33'b1010111001010001_1_1_10_101_001_110_0_x_00;
      patterns[8933] = 33'b1010111001010001_0_0_00_000_000_000_0_0_00;
      patterns[8934] = 33'b1011011001010001_0_1_11_101_001_110_0_x_00;
      patterns[8935] = 33'b1011111001010001_1_1_11_101_001_110_0_x_00;
      patterns[8936] = 33'b1011111001010001_0_0_00_000_000_000_0_0_00;
      patterns[8937] = 33'b0101011001010000_0_1_xx_101_xxx_110_0_1_01;
      patterns[8938] = 33'b0101111001010000_1_1_xx_101_xxx_110_0_1_01;
      patterns[8939] = 33'b0101111001010000_0_0_00_000_000_000_0_0_00;
      patterns[8940] = 33'b0100011001010000_0_0_xx_101_110_xxx_1_x_xx;
      patterns[8941] = 33'b0100111001010000_1_0_xx_101_110_xxx_1_x_xx;
      patterns[8942] = 33'b0100111001010000_0_0_00_000_000_000_0_0_00;
      patterns[8943] = 33'b0000011011000000_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8944] = 33'b0000111011000000_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8945] = 33'b0000111011000000_0_0_00_000_000_000_0_0_00;
      patterns[8946] = 33'b1000011001010010_0_1_00_101_010_110_0_x_00;
      patterns[8947] = 33'b1000111001010010_1_1_00_101_010_110_0_x_00;
      patterns[8948] = 33'b1000111001010010_0_0_00_000_000_000_0_0_00;
      patterns[8949] = 33'b1001011001010010_0_1_01_101_010_110_0_x_00;
      patterns[8950] = 33'b1001111001010010_1_1_01_101_010_110_0_x_00;
      patterns[8951] = 33'b1001111001010010_0_0_00_000_000_000_0_0_00;
      patterns[8952] = 33'b1010011001010010_0_1_10_101_010_110_0_x_00;
      patterns[8953] = 33'b1010111001010010_1_1_10_101_010_110_0_x_00;
      patterns[8954] = 33'b1010111001010010_0_0_00_000_000_000_0_0_00;
      patterns[8955] = 33'b1011011001010010_0_1_11_101_010_110_0_x_00;
      patterns[8956] = 33'b1011111001010010_1_1_11_101_010_110_0_x_00;
      patterns[8957] = 33'b1011111001010010_0_0_00_000_000_000_0_0_00;
      patterns[8958] = 33'b0101011001010000_0_1_xx_101_xxx_110_0_1_01;
      patterns[8959] = 33'b0101111001010000_1_1_xx_101_xxx_110_0_1_01;
      patterns[8960] = 33'b0101111001010000_0_0_00_000_000_000_0_0_00;
      patterns[8961] = 33'b0100011001010000_0_0_xx_101_110_xxx_1_x_xx;
      patterns[8962] = 33'b0100111001010000_1_0_xx_101_110_xxx_1_x_xx;
      patterns[8963] = 33'b0100111001010000_0_0_00_000_000_000_0_0_00;
      patterns[8964] = 33'b0000011001101010_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8965] = 33'b0000111001101010_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8966] = 33'b0000111001101010_0_0_00_000_000_000_0_0_00;
      patterns[8967] = 33'b1000011001010011_0_1_00_101_011_110_0_x_00;
      patterns[8968] = 33'b1000111001010011_1_1_00_101_011_110_0_x_00;
      patterns[8969] = 33'b1000111001010011_0_0_00_000_000_000_0_0_00;
      patterns[8970] = 33'b1001011001010011_0_1_01_101_011_110_0_x_00;
      patterns[8971] = 33'b1001111001010011_1_1_01_101_011_110_0_x_00;
      patterns[8972] = 33'b1001111001010011_0_0_00_000_000_000_0_0_00;
      patterns[8973] = 33'b1010011001010011_0_1_10_101_011_110_0_x_00;
      patterns[8974] = 33'b1010111001010011_1_1_10_101_011_110_0_x_00;
      patterns[8975] = 33'b1010111001010011_0_0_00_000_000_000_0_0_00;
      patterns[8976] = 33'b1011011001010011_0_1_11_101_011_110_0_x_00;
      patterns[8977] = 33'b1011111001010011_1_1_11_101_011_110_0_x_00;
      patterns[8978] = 33'b1011111001010011_0_0_00_000_000_000_0_0_00;
      patterns[8979] = 33'b0101011001010000_0_1_xx_101_xxx_110_0_1_01;
      patterns[8980] = 33'b0101111001010000_1_1_xx_101_xxx_110_0_1_01;
      patterns[8981] = 33'b0101111001010000_0_0_00_000_000_000_0_0_00;
      patterns[8982] = 33'b0100011001010000_0_0_xx_101_110_xxx_1_x_xx;
      patterns[8983] = 33'b0100111001010000_1_0_xx_101_110_xxx_1_x_xx;
      patterns[8984] = 33'b0100111001010000_0_0_00_000_000_000_0_0_00;
      patterns[8985] = 33'b0000011001111111_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[8986] = 33'b0000111001111111_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[8987] = 33'b0000111001111111_0_0_00_000_000_000_0_0_00;
      patterns[8988] = 33'b1000011001010100_0_1_00_101_100_110_0_x_00;
      patterns[8989] = 33'b1000111001010100_1_1_00_101_100_110_0_x_00;
      patterns[8990] = 33'b1000111001010100_0_0_00_000_000_000_0_0_00;
      patterns[8991] = 33'b1001011001010100_0_1_01_101_100_110_0_x_00;
      patterns[8992] = 33'b1001111001010100_1_1_01_101_100_110_0_x_00;
      patterns[8993] = 33'b1001111001010100_0_0_00_000_000_000_0_0_00;
      patterns[8994] = 33'b1010011001010100_0_1_10_101_100_110_0_x_00;
      patterns[8995] = 33'b1010111001010100_1_1_10_101_100_110_0_x_00;
      patterns[8996] = 33'b1010111001010100_0_0_00_000_000_000_0_0_00;
      patterns[8997] = 33'b1011011001010100_0_1_11_101_100_110_0_x_00;
      patterns[8998] = 33'b1011111001010100_1_1_11_101_100_110_0_x_00;
      patterns[8999] = 33'b1011111001010100_0_0_00_000_000_000_0_0_00;
      patterns[9000] = 33'b0101011001010000_0_1_xx_101_xxx_110_0_1_01;
      patterns[9001] = 33'b0101111001010000_1_1_xx_101_xxx_110_0_1_01;
      patterns[9002] = 33'b0101111001010000_0_0_00_000_000_000_0_0_00;
      patterns[9003] = 33'b0100011001010000_0_0_xx_101_110_xxx_1_x_xx;
      patterns[9004] = 33'b0100111001010000_1_0_xx_101_110_xxx_1_x_xx;
      patterns[9005] = 33'b0100111001010000_0_0_00_000_000_000_0_0_00;
      patterns[9006] = 33'b0000011011010111_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9007] = 33'b0000111011010111_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9008] = 33'b0000111011010111_0_0_00_000_000_000_0_0_00;
      patterns[9009] = 33'b1000011001010101_0_1_00_101_101_110_0_x_00;
      patterns[9010] = 33'b1000111001010101_1_1_00_101_101_110_0_x_00;
      patterns[9011] = 33'b1000111001010101_0_0_00_000_000_000_0_0_00;
      patterns[9012] = 33'b1001011001010101_0_1_01_101_101_110_0_x_00;
      patterns[9013] = 33'b1001111001010101_1_1_01_101_101_110_0_x_00;
      patterns[9014] = 33'b1001111001010101_0_0_00_000_000_000_0_0_00;
      patterns[9015] = 33'b1010011001010101_0_1_10_101_101_110_0_x_00;
      patterns[9016] = 33'b1010111001010101_1_1_10_101_101_110_0_x_00;
      patterns[9017] = 33'b1010111001010101_0_0_00_000_000_000_0_0_00;
      patterns[9018] = 33'b1011011001010101_0_1_11_101_101_110_0_x_00;
      patterns[9019] = 33'b1011111001010101_1_1_11_101_101_110_0_x_00;
      patterns[9020] = 33'b1011111001010101_0_0_00_000_000_000_0_0_00;
      patterns[9021] = 33'b0101011001010000_0_1_xx_101_xxx_110_0_1_01;
      patterns[9022] = 33'b0101111001010000_1_1_xx_101_xxx_110_0_1_01;
      patterns[9023] = 33'b0101111001010000_0_0_00_000_000_000_0_0_00;
      patterns[9024] = 33'b0100011001010000_0_0_xx_101_110_xxx_1_x_xx;
      patterns[9025] = 33'b0100111001010000_1_0_xx_101_110_xxx_1_x_xx;
      patterns[9026] = 33'b0100111001010000_0_0_00_000_000_000_0_0_00;
      patterns[9027] = 33'b0000011001011001_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9028] = 33'b0000111001011001_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9029] = 33'b0000111001011001_0_0_00_000_000_000_0_0_00;
      patterns[9030] = 33'b1000011001010110_0_1_00_101_110_110_0_x_00;
      patterns[9031] = 33'b1000111001010110_1_1_00_101_110_110_0_x_00;
      patterns[9032] = 33'b1000111001010110_0_0_00_000_000_000_0_0_00;
      patterns[9033] = 33'b1001011001010110_0_1_01_101_110_110_0_x_00;
      patterns[9034] = 33'b1001111001010110_1_1_01_101_110_110_0_x_00;
      patterns[9035] = 33'b1001111001010110_0_0_00_000_000_000_0_0_00;
      patterns[9036] = 33'b1010011001010110_0_1_10_101_110_110_0_x_00;
      patterns[9037] = 33'b1010111001010110_1_1_10_101_110_110_0_x_00;
      patterns[9038] = 33'b1010111001010110_0_0_00_000_000_000_0_0_00;
      patterns[9039] = 33'b1011011001010110_0_1_11_101_110_110_0_x_00;
      patterns[9040] = 33'b1011111001010110_1_1_11_101_110_110_0_x_00;
      patterns[9041] = 33'b1011111001010110_0_0_00_000_000_000_0_0_00;
      patterns[9042] = 33'b0101011001010000_0_1_xx_101_xxx_110_0_1_01;
      patterns[9043] = 33'b0101111001010000_1_1_xx_101_xxx_110_0_1_01;
      patterns[9044] = 33'b0101111001010000_0_0_00_000_000_000_0_0_00;
      patterns[9045] = 33'b0100011001010000_0_0_xx_101_110_xxx_1_x_xx;
      patterns[9046] = 33'b0100111001010000_1_0_xx_101_110_xxx_1_x_xx;
      patterns[9047] = 33'b0100111001010000_0_0_00_000_000_000_0_0_00;
      patterns[9048] = 33'b0000011001110011_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9049] = 33'b0000111001110011_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9050] = 33'b0000111001110011_0_0_00_000_000_000_0_0_00;
      patterns[9051] = 33'b1000011001010111_0_1_00_101_111_110_0_x_00;
      patterns[9052] = 33'b1000111001010111_1_1_00_101_111_110_0_x_00;
      patterns[9053] = 33'b1000111001010111_0_0_00_000_000_000_0_0_00;
      patterns[9054] = 33'b1001011001010111_0_1_01_101_111_110_0_x_00;
      patterns[9055] = 33'b1001111001010111_1_1_01_101_111_110_0_x_00;
      patterns[9056] = 33'b1001111001010111_0_0_00_000_000_000_0_0_00;
      patterns[9057] = 33'b1010011001010111_0_1_10_101_111_110_0_x_00;
      patterns[9058] = 33'b1010111001010111_1_1_10_101_111_110_0_x_00;
      patterns[9059] = 33'b1010111001010111_0_0_00_000_000_000_0_0_00;
      patterns[9060] = 33'b1011011001010111_0_1_11_101_111_110_0_x_00;
      patterns[9061] = 33'b1011111001010111_1_1_11_101_111_110_0_x_00;
      patterns[9062] = 33'b1011111001010111_0_0_00_000_000_000_0_0_00;
      patterns[9063] = 33'b0101011001010000_0_1_xx_101_xxx_110_0_1_01;
      patterns[9064] = 33'b0101111001010000_1_1_xx_101_xxx_110_0_1_01;
      patterns[9065] = 33'b0101111001010000_0_0_00_000_000_000_0_0_00;
      patterns[9066] = 33'b0100011001010000_0_0_xx_101_110_xxx_1_x_xx;
      patterns[9067] = 33'b0100111001010000_1_0_xx_101_110_xxx_1_x_xx;
      patterns[9068] = 33'b0100111001010000_0_0_00_000_000_000_0_0_00;
      patterns[9069] = 33'b0000011001111010_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9070] = 33'b0000111001111010_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9071] = 33'b0000111001111010_0_0_00_000_000_000_0_0_00;
      patterns[9072] = 33'b1000011001100000_0_1_00_110_000_110_0_x_00;
      patterns[9073] = 33'b1000111001100000_1_1_00_110_000_110_0_x_00;
      patterns[9074] = 33'b1000111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9075] = 33'b1001011001100000_0_1_01_110_000_110_0_x_00;
      patterns[9076] = 33'b1001111001100000_1_1_01_110_000_110_0_x_00;
      patterns[9077] = 33'b1001111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9078] = 33'b1010011001100000_0_1_10_110_000_110_0_x_00;
      patterns[9079] = 33'b1010111001100000_1_1_10_110_000_110_0_x_00;
      patterns[9080] = 33'b1010111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9081] = 33'b1011011001100000_0_1_11_110_000_110_0_x_00;
      patterns[9082] = 33'b1011111001100000_1_1_11_110_000_110_0_x_00;
      patterns[9083] = 33'b1011111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9084] = 33'b0101011001100000_0_1_xx_110_xxx_110_0_1_01;
      patterns[9085] = 33'b0101111001100000_1_1_xx_110_xxx_110_0_1_01;
      patterns[9086] = 33'b0101111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9087] = 33'b0100011001100000_0_0_xx_110_110_xxx_1_x_xx;
      patterns[9088] = 33'b0100111001100000_1_0_xx_110_110_xxx_1_x_xx;
      patterns[9089] = 33'b0100111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9090] = 33'b0000011011101111_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9091] = 33'b0000111011101111_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9092] = 33'b0000111011101111_0_0_00_000_000_000_0_0_00;
      patterns[9093] = 33'b1000011001100001_0_1_00_110_001_110_0_x_00;
      patterns[9094] = 33'b1000111001100001_1_1_00_110_001_110_0_x_00;
      patterns[9095] = 33'b1000111001100001_0_0_00_000_000_000_0_0_00;
      patterns[9096] = 33'b1001011001100001_0_1_01_110_001_110_0_x_00;
      patterns[9097] = 33'b1001111001100001_1_1_01_110_001_110_0_x_00;
      patterns[9098] = 33'b1001111001100001_0_0_00_000_000_000_0_0_00;
      patterns[9099] = 33'b1010011001100001_0_1_10_110_001_110_0_x_00;
      patterns[9100] = 33'b1010111001100001_1_1_10_110_001_110_0_x_00;
      patterns[9101] = 33'b1010111001100001_0_0_00_000_000_000_0_0_00;
      patterns[9102] = 33'b1011011001100001_0_1_11_110_001_110_0_x_00;
      patterns[9103] = 33'b1011111001100001_1_1_11_110_001_110_0_x_00;
      patterns[9104] = 33'b1011111001100001_0_0_00_000_000_000_0_0_00;
      patterns[9105] = 33'b0101011001100000_0_1_xx_110_xxx_110_0_1_01;
      patterns[9106] = 33'b0101111001100000_1_1_xx_110_xxx_110_0_1_01;
      patterns[9107] = 33'b0101111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9108] = 33'b0100011001100000_0_0_xx_110_110_xxx_1_x_xx;
      patterns[9109] = 33'b0100111001100000_1_0_xx_110_110_xxx_1_x_xx;
      patterns[9110] = 33'b0100111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9111] = 33'b0000011010000100_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9112] = 33'b0000111010000100_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9113] = 33'b0000111010000100_0_0_00_000_000_000_0_0_00;
      patterns[9114] = 33'b1000011001100010_0_1_00_110_010_110_0_x_00;
      patterns[9115] = 33'b1000111001100010_1_1_00_110_010_110_0_x_00;
      patterns[9116] = 33'b1000111001100010_0_0_00_000_000_000_0_0_00;
      patterns[9117] = 33'b1001011001100010_0_1_01_110_010_110_0_x_00;
      patterns[9118] = 33'b1001111001100010_1_1_01_110_010_110_0_x_00;
      patterns[9119] = 33'b1001111001100010_0_0_00_000_000_000_0_0_00;
      patterns[9120] = 33'b1010011001100010_0_1_10_110_010_110_0_x_00;
      patterns[9121] = 33'b1010111001100010_1_1_10_110_010_110_0_x_00;
      patterns[9122] = 33'b1010111001100010_0_0_00_000_000_000_0_0_00;
      patterns[9123] = 33'b1011011001100010_0_1_11_110_010_110_0_x_00;
      patterns[9124] = 33'b1011111001100010_1_1_11_110_010_110_0_x_00;
      patterns[9125] = 33'b1011111001100010_0_0_00_000_000_000_0_0_00;
      patterns[9126] = 33'b0101011001100000_0_1_xx_110_xxx_110_0_1_01;
      patterns[9127] = 33'b0101111001100000_1_1_xx_110_xxx_110_0_1_01;
      patterns[9128] = 33'b0101111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9129] = 33'b0100011001100000_0_0_xx_110_110_xxx_1_x_xx;
      patterns[9130] = 33'b0100111001100000_1_0_xx_110_110_xxx_1_x_xx;
      patterns[9131] = 33'b0100111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9132] = 33'b0000011001001001_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9133] = 33'b0000111001001001_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9134] = 33'b0000111001001001_0_0_00_000_000_000_0_0_00;
      patterns[9135] = 33'b1000011001100011_0_1_00_110_011_110_0_x_00;
      patterns[9136] = 33'b1000111001100011_1_1_00_110_011_110_0_x_00;
      patterns[9137] = 33'b1000111001100011_0_0_00_000_000_000_0_0_00;
      patterns[9138] = 33'b1001011001100011_0_1_01_110_011_110_0_x_00;
      patterns[9139] = 33'b1001111001100011_1_1_01_110_011_110_0_x_00;
      patterns[9140] = 33'b1001111001100011_0_0_00_000_000_000_0_0_00;
      patterns[9141] = 33'b1010011001100011_0_1_10_110_011_110_0_x_00;
      patterns[9142] = 33'b1010111001100011_1_1_10_110_011_110_0_x_00;
      patterns[9143] = 33'b1010111001100011_0_0_00_000_000_000_0_0_00;
      patterns[9144] = 33'b1011011001100011_0_1_11_110_011_110_0_x_00;
      patterns[9145] = 33'b1011111001100011_1_1_11_110_011_110_0_x_00;
      patterns[9146] = 33'b1011111001100011_0_0_00_000_000_000_0_0_00;
      patterns[9147] = 33'b0101011001100000_0_1_xx_110_xxx_110_0_1_01;
      patterns[9148] = 33'b0101111001100000_1_1_xx_110_xxx_110_0_1_01;
      patterns[9149] = 33'b0101111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9150] = 33'b0100011001100000_0_0_xx_110_110_xxx_1_x_xx;
      patterns[9151] = 33'b0100111001100000_1_0_xx_110_110_xxx_1_x_xx;
      patterns[9152] = 33'b0100111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9153] = 33'b0000011010000101_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9154] = 33'b0000111010000101_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9155] = 33'b0000111010000101_0_0_00_000_000_000_0_0_00;
      patterns[9156] = 33'b1000011001100100_0_1_00_110_100_110_0_x_00;
      patterns[9157] = 33'b1000111001100100_1_1_00_110_100_110_0_x_00;
      patterns[9158] = 33'b1000111001100100_0_0_00_000_000_000_0_0_00;
      patterns[9159] = 33'b1001011001100100_0_1_01_110_100_110_0_x_00;
      patterns[9160] = 33'b1001111001100100_1_1_01_110_100_110_0_x_00;
      patterns[9161] = 33'b1001111001100100_0_0_00_000_000_000_0_0_00;
      patterns[9162] = 33'b1010011001100100_0_1_10_110_100_110_0_x_00;
      patterns[9163] = 33'b1010111001100100_1_1_10_110_100_110_0_x_00;
      patterns[9164] = 33'b1010111001100100_0_0_00_000_000_000_0_0_00;
      patterns[9165] = 33'b1011011001100100_0_1_11_110_100_110_0_x_00;
      patterns[9166] = 33'b1011111001100100_1_1_11_110_100_110_0_x_00;
      patterns[9167] = 33'b1011111001100100_0_0_00_000_000_000_0_0_00;
      patterns[9168] = 33'b0101011001100000_0_1_xx_110_xxx_110_0_1_01;
      patterns[9169] = 33'b0101111001100000_1_1_xx_110_xxx_110_0_1_01;
      patterns[9170] = 33'b0101111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9171] = 33'b0100011001100000_0_0_xx_110_110_xxx_1_x_xx;
      patterns[9172] = 33'b0100111001100000_1_0_xx_110_110_xxx_1_x_xx;
      patterns[9173] = 33'b0100111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9174] = 33'b0000011000111111_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9175] = 33'b0000111000111111_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9176] = 33'b0000111000111111_0_0_00_000_000_000_0_0_00;
      patterns[9177] = 33'b1000011001100101_0_1_00_110_101_110_0_x_00;
      patterns[9178] = 33'b1000111001100101_1_1_00_110_101_110_0_x_00;
      patterns[9179] = 33'b1000111001100101_0_0_00_000_000_000_0_0_00;
      patterns[9180] = 33'b1001011001100101_0_1_01_110_101_110_0_x_00;
      patterns[9181] = 33'b1001111001100101_1_1_01_110_101_110_0_x_00;
      patterns[9182] = 33'b1001111001100101_0_0_00_000_000_000_0_0_00;
      patterns[9183] = 33'b1010011001100101_0_1_10_110_101_110_0_x_00;
      patterns[9184] = 33'b1010111001100101_1_1_10_110_101_110_0_x_00;
      patterns[9185] = 33'b1010111001100101_0_0_00_000_000_000_0_0_00;
      patterns[9186] = 33'b1011011001100101_0_1_11_110_101_110_0_x_00;
      patterns[9187] = 33'b1011111001100101_1_1_11_110_101_110_0_x_00;
      patterns[9188] = 33'b1011111001100101_0_0_00_000_000_000_0_0_00;
      patterns[9189] = 33'b0101011001100000_0_1_xx_110_xxx_110_0_1_01;
      patterns[9190] = 33'b0101111001100000_1_1_xx_110_xxx_110_0_1_01;
      patterns[9191] = 33'b0101111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9192] = 33'b0100011001100000_0_0_xx_110_110_xxx_1_x_xx;
      patterns[9193] = 33'b0100111001100000_1_0_xx_110_110_xxx_1_x_xx;
      patterns[9194] = 33'b0100111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9195] = 33'b0000011010110111_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9196] = 33'b0000111010110111_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9197] = 33'b0000111010110111_0_0_00_000_000_000_0_0_00;
      patterns[9198] = 33'b1000011001100110_0_1_00_110_110_110_0_x_00;
      patterns[9199] = 33'b1000111001100110_1_1_00_110_110_110_0_x_00;
      patterns[9200] = 33'b1000111001100110_0_0_00_000_000_000_0_0_00;
      patterns[9201] = 33'b1001011001100110_0_1_01_110_110_110_0_x_00;
      patterns[9202] = 33'b1001111001100110_1_1_01_110_110_110_0_x_00;
      patterns[9203] = 33'b1001111001100110_0_0_00_000_000_000_0_0_00;
      patterns[9204] = 33'b1010011001100110_0_1_10_110_110_110_0_x_00;
      patterns[9205] = 33'b1010111001100110_1_1_10_110_110_110_0_x_00;
      patterns[9206] = 33'b1010111001100110_0_0_00_000_000_000_0_0_00;
      patterns[9207] = 33'b1011011001100110_0_1_11_110_110_110_0_x_00;
      patterns[9208] = 33'b1011111001100110_1_1_11_110_110_110_0_x_00;
      patterns[9209] = 33'b1011111001100110_0_0_00_000_000_000_0_0_00;
      patterns[9210] = 33'b0101011001100000_0_1_xx_110_xxx_110_0_1_01;
      patterns[9211] = 33'b0101111001100000_1_1_xx_110_xxx_110_0_1_01;
      patterns[9212] = 33'b0101111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9213] = 33'b0100011001100000_0_0_xx_110_110_xxx_1_x_xx;
      patterns[9214] = 33'b0100111001100000_1_0_xx_110_110_xxx_1_x_xx;
      patterns[9215] = 33'b0100111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9216] = 33'b0000011010001001_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9217] = 33'b0000111010001001_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9218] = 33'b0000111010001001_0_0_00_000_000_000_0_0_00;
      patterns[9219] = 33'b1000011001100111_0_1_00_110_111_110_0_x_00;
      patterns[9220] = 33'b1000111001100111_1_1_00_110_111_110_0_x_00;
      patterns[9221] = 33'b1000111001100111_0_0_00_000_000_000_0_0_00;
      patterns[9222] = 33'b1001011001100111_0_1_01_110_111_110_0_x_00;
      patterns[9223] = 33'b1001111001100111_1_1_01_110_111_110_0_x_00;
      patterns[9224] = 33'b1001111001100111_0_0_00_000_000_000_0_0_00;
      patterns[9225] = 33'b1010011001100111_0_1_10_110_111_110_0_x_00;
      patterns[9226] = 33'b1010111001100111_1_1_10_110_111_110_0_x_00;
      patterns[9227] = 33'b1010111001100111_0_0_00_000_000_000_0_0_00;
      patterns[9228] = 33'b1011011001100111_0_1_11_110_111_110_0_x_00;
      patterns[9229] = 33'b1011111001100111_1_1_11_110_111_110_0_x_00;
      patterns[9230] = 33'b1011111001100111_0_0_00_000_000_000_0_0_00;
      patterns[9231] = 33'b0101011001100000_0_1_xx_110_xxx_110_0_1_01;
      patterns[9232] = 33'b0101111001100000_1_1_xx_110_xxx_110_0_1_01;
      patterns[9233] = 33'b0101111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9234] = 33'b0100011001100000_0_0_xx_110_110_xxx_1_x_xx;
      patterns[9235] = 33'b0100111001100000_1_0_xx_110_110_xxx_1_x_xx;
      patterns[9236] = 33'b0100111001100000_0_0_00_000_000_000_0_0_00;
      patterns[9237] = 33'b0000011011111000_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9238] = 33'b0000111011111000_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9239] = 33'b0000111011111000_0_0_00_000_000_000_0_0_00;
      patterns[9240] = 33'b1000011001110000_0_1_00_111_000_110_0_x_00;
      patterns[9241] = 33'b1000111001110000_1_1_00_111_000_110_0_x_00;
      patterns[9242] = 33'b1000111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9243] = 33'b1001011001110000_0_1_01_111_000_110_0_x_00;
      patterns[9244] = 33'b1001111001110000_1_1_01_111_000_110_0_x_00;
      patterns[9245] = 33'b1001111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9246] = 33'b1010011001110000_0_1_10_111_000_110_0_x_00;
      patterns[9247] = 33'b1010111001110000_1_1_10_111_000_110_0_x_00;
      patterns[9248] = 33'b1010111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9249] = 33'b1011011001110000_0_1_11_111_000_110_0_x_00;
      patterns[9250] = 33'b1011111001110000_1_1_11_111_000_110_0_x_00;
      patterns[9251] = 33'b1011111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9252] = 33'b0101011001110000_0_1_xx_111_xxx_110_0_1_01;
      patterns[9253] = 33'b0101111001110000_1_1_xx_111_xxx_110_0_1_01;
      patterns[9254] = 33'b0101111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9255] = 33'b0100011001110000_0_0_xx_111_110_xxx_1_x_xx;
      patterns[9256] = 33'b0100111001110000_1_0_xx_111_110_xxx_1_x_xx;
      patterns[9257] = 33'b0100111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9258] = 33'b0000011001101110_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9259] = 33'b0000111001101110_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9260] = 33'b0000111001101110_0_0_00_000_000_000_0_0_00;
      patterns[9261] = 33'b1000011001110001_0_1_00_111_001_110_0_x_00;
      patterns[9262] = 33'b1000111001110001_1_1_00_111_001_110_0_x_00;
      patterns[9263] = 33'b1000111001110001_0_0_00_000_000_000_0_0_00;
      patterns[9264] = 33'b1001011001110001_0_1_01_111_001_110_0_x_00;
      patterns[9265] = 33'b1001111001110001_1_1_01_111_001_110_0_x_00;
      patterns[9266] = 33'b1001111001110001_0_0_00_000_000_000_0_0_00;
      patterns[9267] = 33'b1010011001110001_0_1_10_111_001_110_0_x_00;
      patterns[9268] = 33'b1010111001110001_1_1_10_111_001_110_0_x_00;
      patterns[9269] = 33'b1010111001110001_0_0_00_000_000_000_0_0_00;
      patterns[9270] = 33'b1011011001110001_0_1_11_111_001_110_0_x_00;
      patterns[9271] = 33'b1011111001110001_1_1_11_111_001_110_0_x_00;
      patterns[9272] = 33'b1011111001110001_0_0_00_000_000_000_0_0_00;
      patterns[9273] = 33'b0101011001110000_0_1_xx_111_xxx_110_0_1_01;
      patterns[9274] = 33'b0101111001110000_1_1_xx_111_xxx_110_0_1_01;
      patterns[9275] = 33'b0101111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9276] = 33'b0100011001110000_0_0_xx_111_110_xxx_1_x_xx;
      patterns[9277] = 33'b0100111001110000_1_0_xx_111_110_xxx_1_x_xx;
      patterns[9278] = 33'b0100111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9279] = 33'b0000011001011101_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9280] = 33'b0000111001011101_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9281] = 33'b0000111001011101_0_0_00_000_000_000_0_0_00;
      patterns[9282] = 33'b1000011001110010_0_1_00_111_010_110_0_x_00;
      patterns[9283] = 33'b1000111001110010_1_1_00_111_010_110_0_x_00;
      patterns[9284] = 33'b1000111001110010_0_0_00_000_000_000_0_0_00;
      patterns[9285] = 33'b1001011001110010_0_1_01_111_010_110_0_x_00;
      patterns[9286] = 33'b1001111001110010_1_1_01_111_010_110_0_x_00;
      patterns[9287] = 33'b1001111001110010_0_0_00_000_000_000_0_0_00;
      patterns[9288] = 33'b1010011001110010_0_1_10_111_010_110_0_x_00;
      patterns[9289] = 33'b1010111001110010_1_1_10_111_010_110_0_x_00;
      patterns[9290] = 33'b1010111001110010_0_0_00_000_000_000_0_0_00;
      patterns[9291] = 33'b1011011001110010_0_1_11_111_010_110_0_x_00;
      patterns[9292] = 33'b1011111001110010_1_1_11_111_010_110_0_x_00;
      patterns[9293] = 33'b1011111001110010_0_0_00_000_000_000_0_0_00;
      patterns[9294] = 33'b0101011001110000_0_1_xx_111_xxx_110_0_1_01;
      patterns[9295] = 33'b0101111001110000_1_1_xx_111_xxx_110_0_1_01;
      patterns[9296] = 33'b0101111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9297] = 33'b0100011001110000_0_0_xx_111_110_xxx_1_x_xx;
      patterns[9298] = 33'b0100111001110000_1_0_xx_111_110_xxx_1_x_xx;
      patterns[9299] = 33'b0100111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9300] = 33'b0000011010111101_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9301] = 33'b0000111010111101_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9302] = 33'b0000111010111101_0_0_00_000_000_000_0_0_00;
      patterns[9303] = 33'b1000011001110011_0_1_00_111_011_110_0_x_00;
      patterns[9304] = 33'b1000111001110011_1_1_00_111_011_110_0_x_00;
      patterns[9305] = 33'b1000111001110011_0_0_00_000_000_000_0_0_00;
      patterns[9306] = 33'b1001011001110011_0_1_01_111_011_110_0_x_00;
      patterns[9307] = 33'b1001111001110011_1_1_01_111_011_110_0_x_00;
      patterns[9308] = 33'b1001111001110011_0_0_00_000_000_000_0_0_00;
      patterns[9309] = 33'b1010011001110011_0_1_10_111_011_110_0_x_00;
      patterns[9310] = 33'b1010111001110011_1_1_10_111_011_110_0_x_00;
      patterns[9311] = 33'b1010111001110011_0_0_00_000_000_000_0_0_00;
      patterns[9312] = 33'b1011011001110011_0_1_11_111_011_110_0_x_00;
      patterns[9313] = 33'b1011111001110011_1_1_11_111_011_110_0_x_00;
      patterns[9314] = 33'b1011111001110011_0_0_00_000_000_000_0_0_00;
      patterns[9315] = 33'b0101011001110000_0_1_xx_111_xxx_110_0_1_01;
      patterns[9316] = 33'b0101111001110000_1_1_xx_111_xxx_110_0_1_01;
      patterns[9317] = 33'b0101111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9318] = 33'b0100011001110000_0_0_xx_111_110_xxx_1_x_xx;
      patterns[9319] = 33'b0100111001110000_1_0_xx_111_110_xxx_1_x_xx;
      patterns[9320] = 33'b0100111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9321] = 33'b0000011011001010_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9322] = 33'b0000111011001010_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9323] = 33'b0000111011001010_0_0_00_000_000_000_0_0_00;
      patterns[9324] = 33'b1000011001110100_0_1_00_111_100_110_0_x_00;
      patterns[9325] = 33'b1000111001110100_1_1_00_111_100_110_0_x_00;
      patterns[9326] = 33'b1000111001110100_0_0_00_000_000_000_0_0_00;
      patterns[9327] = 33'b1001011001110100_0_1_01_111_100_110_0_x_00;
      patterns[9328] = 33'b1001111001110100_1_1_01_111_100_110_0_x_00;
      patterns[9329] = 33'b1001111001110100_0_0_00_000_000_000_0_0_00;
      patterns[9330] = 33'b1010011001110100_0_1_10_111_100_110_0_x_00;
      patterns[9331] = 33'b1010111001110100_1_1_10_111_100_110_0_x_00;
      patterns[9332] = 33'b1010111001110100_0_0_00_000_000_000_0_0_00;
      patterns[9333] = 33'b1011011001110100_0_1_11_111_100_110_0_x_00;
      patterns[9334] = 33'b1011111001110100_1_1_11_111_100_110_0_x_00;
      patterns[9335] = 33'b1011111001110100_0_0_00_000_000_000_0_0_00;
      patterns[9336] = 33'b0101011001110000_0_1_xx_111_xxx_110_0_1_01;
      patterns[9337] = 33'b0101111001110000_1_1_xx_111_xxx_110_0_1_01;
      patterns[9338] = 33'b0101111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9339] = 33'b0100011001110000_0_0_xx_111_110_xxx_1_x_xx;
      patterns[9340] = 33'b0100111001110000_1_0_xx_111_110_xxx_1_x_xx;
      patterns[9341] = 33'b0100111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9342] = 33'b0000011011100010_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9343] = 33'b0000111011100010_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9344] = 33'b0000111011100010_0_0_00_000_000_000_0_0_00;
      patterns[9345] = 33'b1000011001110101_0_1_00_111_101_110_0_x_00;
      patterns[9346] = 33'b1000111001110101_1_1_00_111_101_110_0_x_00;
      patterns[9347] = 33'b1000111001110101_0_0_00_000_000_000_0_0_00;
      patterns[9348] = 33'b1001011001110101_0_1_01_111_101_110_0_x_00;
      patterns[9349] = 33'b1001111001110101_1_1_01_111_101_110_0_x_00;
      patterns[9350] = 33'b1001111001110101_0_0_00_000_000_000_0_0_00;
      patterns[9351] = 33'b1010011001110101_0_1_10_111_101_110_0_x_00;
      patterns[9352] = 33'b1010111001110101_1_1_10_111_101_110_0_x_00;
      patterns[9353] = 33'b1010111001110101_0_0_00_000_000_000_0_0_00;
      patterns[9354] = 33'b1011011001110101_0_1_11_111_101_110_0_x_00;
      patterns[9355] = 33'b1011111001110101_1_1_11_111_101_110_0_x_00;
      patterns[9356] = 33'b1011111001110101_0_0_00_000_000_000_0_0_00;
      patterns[9357] = 33'b0101011001110000_0_1_xx_111_xxx_110_0_1_01;
      patterns[9358] = 33'b0101111001110000_1_1_xx_111_xxx_110_0_1_01;
      patterns[9359] = 33'b0101111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9360] = 33'b0100011001110000_0_0_xx_111_110_xxx_1_x_xx;
      patterns[9361] = 33'b0100111001110000_1_0_xx_111_110_xxx_1_x_xx;
      patterns[9362] = 33'b0100111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9363] = 33'b0000011010111111_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9364] = 33'b0000111010111111_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9365] = 33'b0000111010111111_0_0_00_000_000_000_0_0_00;
      patterns[9366] = 33'b1000011001110110_0_1_00_111_110_110_0_x_00;
      patterns[9367] = 33'b1000111001110110_1_1_00_111_110_110_0_x_00;
      patterns[9368] = 33'b1000111001110110_0_0_00_000_000_000_0_0_00;
      patterns[9369] = 33'b1001011001110110_0_1_01_111_110_110_0_x_00;
      patterns[9370] = 33'b1001111001110110_1_1_01_111_110_110_0_x_00;
      patterns[9371] = 33'b1001111001110110_0_0_00_000_000_000_0_0_00;
      patterns[9372] = 33'b1010011001110110_0_1_10_111_110_110_0_x_00;
      patterns[9373] = 33'b1010111001110110_1_1_10_111_110_110_0_x_00;
      patterns[9374] = 33'b1010111001110110_0_0_00_000_000_000_0_0_00;
      patterns[9375] = 33'b1011011001110110_0_1_11_111_110_110_0_x_00;
      patterns[9376] = 33'b1011111001110110_1_1_11_111_110_110_0_x_00;
      patterns[9377] = 33'b1011111001110110_0_0_00_000_000_000_0_0_00;
      patterns[9378] = 33'b0101011001110000_0_1_xx_111_xxx_110_0_1_01;
      patterns[9379] = 33'b0101111001110000_1_1_xx_111_xxx_110_0_1_01;
      patterns[9380] = 33'b0101111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9381] = 33'b0100011001110000_0_0_xx_111_110_xxx_1_x_xx;
      patterns[9382] = 33'b0100111001110000_1_0_xx_111_110_xxx_1_x_xx;
      patterns[9383] = 33'b0100111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9384] = 33'b0000011000001110_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9385] = 33'b0000111000001110_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9386] = 33'b0000111000001110_0_0_00_000_000_000_0_0_00;
      patterns[9387] = 33'b1000011001110111_0_1_00_111_111_110_0_x_00;
      patterns[9388] = 33'b1000111001110111_1_1_00_111_111_110_0_x_00;
      patterns[9389] = 33'b1000111001110111_0_0_00_000_000_000_0_0_00;
      patterns[9390] = 33'b1001011001110111_0_1_01_111_111_110_0_x_00;
      patterns[9391] = 33'b1001111001110111_1_1_01_111_111_110_0_x_00;
      patterns[9392] = 33'b1001111001110111_0_0_00_000_000_000_0_0_00;
      patterns[9393] = 33'b1010011001110111_0_1_10_111_111_110_0_x_00;
      patterns[9394] = 33'b1010111001110111_1_1_10_111_111_110_0_x_00;
      patterns[9395] = 33'b1010111001110111_0_0_00_000_000_000_0_0_00;
      patterns[9396] = 33'b1011011001110111_0_1_11_111_111_110_0_x_00;
      patterns[9397] = 33'b1011111001110111_1_1_11_111_111_110_0_x_00;
      patterns[9398] = 33'b1011111001110111_0_0_00_000_000_000_0_0_00;
      patterns[9399] = 33'b0101011001110000_0_1_xx_111_xxx_110_0_1_01;
      patterns[9400] = 33'b0101111001110000_1_1_xx_111_xxx_110_0_1_01;
      patterns[9401] = 33'b0101111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9402] = 33'b0100011001110000_0_0_xx_111_110_xxx_1_x_xx;
      patterns[9403] = 33'b0100111001110000_1_0_xx_111_110_xxx_1_x_xx;
      patterns[9404] = 33'b0100111001110000_0_0_00_000_000_000_0_0_00;
      patterns[9405] = 33'b0000011010010000_0_1_xx_xxx_xxx_110_0_x_10;
      patterns[9406] = 33'b0000111010010000_1_1_xx_xxx_xxx_110_0_x_10;
      patterns[9407] = 33'b0000111010010000_0_0_00_000_000_000_0_0_00;
      patterns[9408] = 33'b1000011100000000_0_1_00_000_000_111_0_x_00;
      patterns[9409] = 33'b1000111100000000_1_1_00_000_000_111_0_x_00;
      patterns[9410] = 33'b1000111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9411] = 33'b1001011100000000_0_1_01_000_000_111_0_x_00;
      patterns[9412] = 33'b1001111100000000_1_1_01_000_000_111_0_x_00;
      patterns[9413] = 33'b1001111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9414] = 33'b1010011100000000_0_1_10_000_000_111_0_x_00;
      patterns[9415] = 33'b1010111100000000_1_1_10_000_000_111_0_x_00;
      patterns[9416] = 33'b1010111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9417] = 33'b1011011100000000_0_1_11_000_000_111_0_x_00;
      patterns[9418] = 33'b1011111100000000_1_1_11_000_000_111_0_x_00;
      patterns[9419] = 33'b1011111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9420] = 33'b0101011100000000_0_1_xx_000_xxx_111_0_1_01;
      patterns[9421] = 33'b0101111100000000_1_1_xx_000_xxx_111_0_1_01;
      patterns[9422] = 33'b0101111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9423] = 33'b0100011100000000_0_0_xx_000_111_xxx_1_x_xx;
      patterns[9424] = 33'b0100111100000000_1_0_xx_000_111_xxx_1_x_xx;
      patterns[9425] = 33'b0100111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9426] = 33'b0000011100011110_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9427] = 33'b0000111100011110_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9428] = 33'b0000111100011110_0_0_00_000_000_000_0_0_00;
      patterns[9429] = 33'b1000011100000001_0_1_00_000_001_111_0_x_00;
      patterns[9430] = 33'b1000111100000001_1_1_00_000_001_111_0_x_00;
      patterns[9431] = 33'b1000111100000001_0_0_00_000_000_000_0_0_00;
      patterns[9432] = 33'b1001011100000001_0_1_01_000_001_111_0_x_00;
      patterns[9433] = 33'b1001111100000001_1_1_01_000_001_111_0_x_00;
      patterns[9434] = 33'b1001111100000001_0_0_00_000_000_000_0_0_00;
      patterns[9435] = 33'b1010011100000001_0_1_10_000_001_111_0_x_00;
      patterns[9436] = 33'b1010111100000001_1_1_10_000_001_111_0_x_00;
      patterns[9437] = 33'b1010111100000001_0_0_00_000_000_000_0_0_00;
      patterns[9438] = 33'b1011011100000001_0_1_11_000_001_111_0_x_00;
      patterns[9439] = 33'b1011111100000001_1_1_11_000_001_111_0_x_00;
      patterns[9440] = 33'b1011111100000001_0_0_00_000_000_000_0_0_00;
      patterns[9441] = 33'b0101011100000000_0_1_xx_000_xxx_111_0_1_01;
      patterns[9442] = 33'b0101111100000000_1_1_xx_000_xxx_111_0_1_01;
      patterns[9443] = 33'b0101111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9444] = 33'b0100011100000000_0_0_xx_000_111_xxx_1_x_xx;
      patterns[9445] = 33'b0100111100000000_1_0_xx_000_111_xxx_1_x_xx;
      patterns[9446] = 33'b0100111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9447] = 33'b0000011110111100_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9448] = 33'b0000111110111100_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9449] = 33'b0000111110111100_0_0_00_000_000_000_0_0_00;
      patterns[9450] = 33'b1000011100000010_0_1_00_000_010_111_0_x_00;
      patterns[9451] = 33'b1000111100000010_1_1_00_000_010_111_0_x_00;
      patterns[9452] = 33'b1000111100000010_0_0_00_000_000_000_0_0_00;
      patterns[9453] = 33'b1001011100000010_0_1_01_000_010_111_0_x_00;
      patterns[9454] = 33'b1001111100000010_1_1_01_000_010_111_0_x_00;
      patterns[9455] = 33'b1001111100000010_0_0_00_000_000_000_0_0_00;
      patterns[9456] = 33'b1010011100000010_0_1_10_000_010_111_0_x_00;
      patterns[9457] = 33'b1010111100000010_1_1_10_000_010_111_0_x_00;
      patterns[9458] = 33'b1010111100000010_0_0_00_000_000_000_0_0_00;
      patterns[9459] = 33'b1011011100000010_0_1_11_000_010_111_0_x_00;
      patterns[9460] = 33'b1011111100000010_1_1_11_000_010_111_0_x_00;
      patterns[9461] = 33'b1011111100000010_0_0_00_000_000_000_0_0_00;
      patterns[9462] = 33'b0101011100000000_0_1_xx_000_xxx_111_0_1_01;
      patterns[9463] = 33'b0101111100000000_1_1_xx_000_xxx_111_0_1_01;
      patterns[9464] = 33'b0101111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9465] = 33'b0100011100000000_0_0_xx_000_111_xxx_1_x_xx;
      patterns[9466] = 33'b0100111100000000_1_0_xx_000_111_xxx_1_x_xx;
      patterns[9467] = 33'b0100111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9468] = 33'b0000011111110000_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9469] = 33'b0000111111110000_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9470] = 33'b0000111111110000_0_0_00_000_000_000_0_0_00;
      patterns[9471] = 33'b1000011100000011_0_1_00_000_011_111_0_x_00;
      patterns[9472] = 33'b1000111100000011_1_1_00_000_011_111_0_x_00;
      patterns[9473] = 33'b1000111100000011_0_0_00_000_000_000_0_0_00;
      patterns[9474] = 33'b1001011100000011_0_1_01_000_011_111_0_x_00;
      patterns[9475] = 33'b1001111100000011_1_1_01_000_011_111_0_x_00;
      patterns[9476] = 33'b1001111100000011_0_0_00_000_000_000_0_0_00;
      patterns[9477] = 33'b1010011100000011_0_1_10_000_011_111_0_x_00;
      patterns[9478] = 33'b1010111100000011_1_1_10_000_011_111_0_x_00;
      patterns[9479] = 33'b1010111100000011_0_0_00_000_000_000_0_0_00;
      patterns[9480] = 33'b1011011100000011_0_1_11_000_011_111_0_x_00;
      patterns[9481] = 33'b1011111100000011_1_1_11_000_011_111_0_x_00;
      patterns[9482] = 33'b1011111100000011_0_0_00_000_000_000_0_0_00;
      patterns[9483] = 33'b0101011100000000_0_1_xx_000_xxx_111_0_1_01;
      patterns[9484] = 33'b0101111100000000_1_1_xx_000_xxx_111_0_1_01;
      patterns[9485] = 33'b0101111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9486] = 33'b0100011100000000_0_0_xx_000_111_xxx_1_x_xx;
      patterns[9487] = 33'b0100111100000000_1_0_xx_000_111_xxx_1_x_xx;
      patterns[9488] = 33'b0100111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9489] = 33'b0000011111001101_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9490] = 33'b0000111111001101_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9491] = 33'b0000111111001101_0_0_00_000_000_000_0_0_00;
      patterns[9492] = 33'b1000011100000100_0_1_00_000_100_111_0_x_00;
      patterns[9493] = 33'b1000111100000100_1_1_00_000_100_111_0_x_00;
      patterns[9494] = 33'b1000111100000100_0_0_00_000_000_000_0_0_00;
      patterns[9495] = 33'b1001011100000100_0_1_01_000_100_111_0_x_00;
      patterns[9496] = 33'b1001111100000100_1_1_01_000_100_111_0_x_00;
      patterns[9497] = 33'b1001111100000100_0_0_00_000_000_000_0_0_00;
      patterns[9498] = 33'b1010011100000100_0_1_10_000_100_111_0_x_00;
      patterns[9499] = 33'b1010111100000100_1_1_10_000_100_111_0_x_00;
      patterns[9500] = 33'b1010111100000100_0_0_00_000_000_000_0_0_00;
      patterns[9501] = 33'b1011011100000100_0_1_11_000_100_111_0_x_00;
      patterns[9502] = 33'b1011111100000100_1_1_11_000_100_111_0_x_00;
      patterns[9503] = 33'b1011111100000100_0_0_00_000_000_000_0_0_00;
      patterns[9504] = 33'b0101011100000000_0_1_xx_000_xxx_111_0_1_01;
      patterns[9505] = 33'b0101111100000000_1_1_xx_000_xxx_111_0_1_01;
      patterns[9506] = 33'b0101111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9507] = 33'b0100011100000000_0_0_xx_000_111_xxx_1_x_xx;
      patterns[9508] = 33'b0100111100000000_1_0_xx_000_111_xxx_1_x_xx;
      patterns[9509] = 33'b0100111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9510] = 33'b0000011111110010_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9511] = 33'b0000111111110010_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9512] = 33'b0000111111110010_0_0_00_000_000_000_0_0_00;
      patterns[9513] = 33'b1000011100000101_0_1_00_000_101_111_0_x_00;
      patterns[9514] = 33'b1000111100000101_1_1_00_000_101_111_0_x_00;
      patterns[9515] = 33'b1000111100000101_0_0_00_000_000_000_0_0_00;
      patterns[9516] = 33'b1001011100000101_0_1_01_000_101_111_0_x_00;
      patterns[9517] = 33'b1001111100000101_1_1_01_000_101_111_0_x_00;
      patterns[9518] = 33'b1001111100000101_0_0_00_000_000_000_0_0_00;
      patterns[9519] = 33'b1010011100000101_0_1_10_000_101_111_0_x_00;
      patterns[9520] = 33'b1010111100000101_1_1_10_000_101_111_0_x_00;
      patterns[9521] = 33'b1010111100000101_0_0_00_000_000_000_0_0_00;
      patterns[9522] = 33'b1011011100000101_0_1_11_000_101_111_0_x_00;
      patterns[9523] = 33'b1011111100000101_1_1_11_000_101_111_0_x_00;
      patterns[9524] = 33'b1011111100000101_0_0_00_000_000_000_0_0_00;
      patterns[9525] = 33'b0101011100000000_0_1_xx_000_xxx_111_0_1_01;
      patterns[9526] = 33'b0101111100000000_1_1_xx_000_xxx_111_0_1_01;
      patterns[9527] = 33'b0101111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9528] = 33'b0100011100000000_0_0_xx_000_111_xxx_1_x_xx;
      patterns[9529] = 33'b0100111100000000_1_0_xx_000_111_xxx_1_x_xx;
      patterns[9530] = 33'b0100111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9531] = 33'b0000011100100010_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9532] = 33'b0000111100100010_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9533] = 33'b0000111100100010_0_0_00_000_000_000_0_0_00;
      patterns[9534] = 33'b1000011100000110_0_1_00_000_110_111_0_x_00;
      patterns[9535] = 33'b1000111100000110_1_1_00_000_110_111_0_x_00;
      patterns[9536] = 33'b1000111100000110_0_0_00_000_000_000_0_0_00;
      patterns[9537] = 33'b1001011100000110_0_1_01_000_110_111_0_x_00;
      patterns[9538] = 33'b1001111100000110_1_1_01_000_110_111_0_x_00;
      patterns[9539] = 33'b1001111100000110_0_0_00_000_000_000_0_0_00;
      patterns[9540] = 33'b1010011100000110_0_1_10_000_110_111_0_x_00;
      patterns[9541] = 33'b1010111100000110_1_1_10_000_110_111_0_x_00;
      patterns[9542] = 33'b1010111100000110_0_0_00_000_000_000_0_0_00;
      patterns[9543] = 33'b1011011100000110_0_1_11_000_110_111_0_x_00;
      patterns[9544] = 33'b1011111100000110_1_1_11_000_110_111_0_x_00;
      patterns[9545] = 33'b1011111100000110_0_0_00_000_000_000_0_0_00;
      patterns[9546] = 33'b0101011100000000_0_1_xx_000_xxx_111_0_1_01;
      patterns[9547] = 33'b0101111100000000_1_1_xx_000_xxx_111_0_1_01;
      patterns[9548] = 33'b0101111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9549] = 33'b0100011100000000_0_0_xx_000_111_xxx_1_x_xx;
      patterns[9550] = 33'b0100111100000000_1_0_xx_000_111_xxx_1_x_xx;
      patterns[9551] = 33'b0100111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9552] = 33'b0000011101101101_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9553] = 33'b0000111101101101_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9554] = 33'b0000111101101101_0_0_00_000_000_000_0_0_00;
      patterns[9555] = 33'b1000011100000111_0_1_00_000_111_111_0_x_00;
      patterns[9556] = 33'b1000111100000111_1_1_00_000_111_111_0_x_00;
      patterns[9557] = 33'b1000111100000111_0_0_00_000_000_000_0_0_00;
      patterns[9558] = 33'b1001011100000111_0_1_01_000_111_111_0_x_00;
      patterns[9559] = 33'b1001111100000111_1_1_01_000_111_111_0_x_00;
      patterns[9560] = 33'b1001111100000111_0_0_00_000_000_000_0_0_00;
      patterns[9561] = 33'b1010011100000111_0_1_10_000_111_111_0_x_00;
      patterns[9562] = 33'b1010111100000111_1_1_10_000_111_111_0_x_00;
      patterns[9563] = 33'b1010111100000111_0_0_00_000_000_000_0_0_00;
      patterns[9564] = 33'b1011011100000111_0_1_11_000_111_111_0_x_00;
      patterns[9565] = 33'b1011111100000111_1_1_11_000_111_111_0_x_00;
      patterns[9566] = 33'b1011111100000111_0_0_00_000_000_000_0_0_00;
      patterns[9567] = 33'b0101011100000000_0_1_xx_000_xxx_111_0_1_01;
      patterns[9568] = 33'b0101111100000000_1_1_xx_000_xxx_111_0_1_01;
      patterns[9569] = 33'b0101111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9570] = 33'b0100011100000000_0_0_xx_000_111_xxx_1_x_xx;
      patterns[9571] = 33'b0100111100000000_1_0_xx_000_111_xxx_1_x_xx;
      patterns[9572] = 33'b0100111100000000_0_0_00_000_000_000_0_0_00;
      patterns[9573] = 33'b0000011110101111_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9574] = 33'b0000111110101111_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9575] = 33'b0000111110101111_0_0_00_000_000_000_0_0_00;
      patterns[9576] = 33'b1000011100010000_0_1_00_001_000_111_0_x_00;
      patterns[9577] = 33'b1000111100010000_1_1_00_001_000_111_0_x_00;
      patterns[9578] = 33'b1000111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9579] = 33'b1001011100010000_0_1_01_001_000_111_0_x_00;
      patterns[9580] = 33'b1001111100010000_1_1_01_001_000_111_0_x_00;
      patterns[9581] = 33'b1001111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9582] = 33'b1010011100010000_0_1_10_001_000_111_0_x_00;
      patterns[9583] = 33'b1010111100010000_1_1_10_001_000_111_0_x_00;
      patterns[9584] = 33'b1010111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9585] = 33'b1011011100010000_0_1_11_001_000_111_0_x_00;
      patterns[9586] = 33'b1011111100010000_1_1_11_001_000_111_0_x_00;
      patterns[9587] = 33'b1011111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9588] = 33'b0101011100010000_0_1_xx_001_xxx_111_0_1_01;
      patterns[9589] = 33'b0101111100010000_1_1_xx_001_xxx_111_0_1_01;
      patterns[9590] = 33'b0101111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9591] = 33'b0100011100010000_0_0_xx_001_111_xxx_1_x_xx;
      patterns[9592] = 33'b0100111100010000_1_0_xx_001_111_xxx_1_x_xx;
      patterns[9593] = 33'b0100111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9594] = 33'b0000011111100110_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9595] = 33'b0000111111100110_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9596] = 33'b0000111111100110_0_0_00_000_000_000_0_0_00;
      patterns[9597] = 33'b1000011100010001_0_1_00_001_001_111_0_x_00;
      patterns[9598] = 33'b1000111100010001_1_1_00_001_001_111_0_x_00;
      patterns[9599] = 33'b1000111100010001_0_0_00_000_000_000_0_0_00;
      patterns[9600] = 33'b1001011100010001_0_1_01_001_001_111_0_x_00;
      patterns[9601] = 33'b1001111100010001_1_1_01_001_001_111_0_x_00;
      patterns[9602] = 33'b1001111100010001_0_0_00_000_000_000_0_0_00;
      patterns[9603] = 33'b1010011100010001_0_1_10_001_001_111_0_x_00;
      patterns[9604] = 33'b1010111100010001_1_1_10_001_001_111_0_x_00;
      patterns[9605] = 33'b1010111100010001_0_0_00_000_000_000_0_0_00;
      patterns[9606] = 33'b1011011100010001_0_1_11_001_001_111_0_x_00;
      patterns[9607] = 33'b1011111100010001_1_1_11_001_001_111_0_x_00;
      patterns[9608] = 33'b1011111100010001_0_0_00_000_000_000_0_0_00;
      patterns[9609] = 33'b0101011100010000_0_1_xx_001_xxx_111_0_1_01;
      patterns[9610] = 33'b0101111100010000_1_1_xx_001_xxx_111_0_1_01;
      patterns[9611] = 33'b0101111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9612] = 33'b0100011100010000_0_0_xx_001_111_xxx_1_x_xx;
      patterns[9613] = 33'b0100111100010000_1_0_xx_001_111_xxx_1_x_xx;
      patterns[9614] = 33'b0100111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9615] = 33'b0000011111010101_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9616] = 33'b0000111111010101_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9617] = 33'b0000111111010101_0_0_00_000_000_000_0_0_00;
      patterns[9618] = 33'b1000011100010010_0_1_00_001_010_111_0_x_00;
      patterns[9619] = 33'b1000111100010010_1_1_00_001_010_111_0_x_00;
      patterns[9620] = 33'b1000111100010010_0_0_00_000_000_000_0_0_00;
      patterns[9621] = 33'b1001011100010010_0_1_01_001_010_111_0_x_00;
      patterns[9622] = 33'b1001111100010010_1_1_01_001_010_111_0_x_00;
      patterns[9623] = 33'b1001111100010010_0_0_00_000_000_000_0_0_00;
      patterns[9624] = 33'b1010011100010010_0_1_10_001_010_111_0_x_00;
      patterns[9625] = 33'b1010111100010010_1_1_10_001_010_111_0_x_00;
      patterns[9626] = 33'b1010111100010010_0_0_00_000_000_000_0_0_00;
      patterns[9627] = 33'b1011011100010010_0_1_11_001_010_111_0_x_00;
      patterns[9628] = 33'b1011111100010010_1_1_11_001_010_111_0_x_00;
      patterns[9629] = 33'b1011111100010010_0_0_00_000_000_000_0_0_00;
      patterns[9630] = 33'b0101011100010000_0_1_xx_001_xxx_111_0_1_01;
      patterns[9631] = 33'b0101111100010000_1_1_xx_001_xxx_111_0_1_01;
      patterns[9632] = 33'b0101111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9633] = 33'b0100011100010000_0_0_xx_001_111_xxx_1_x_xx;
      patterns[9634] = 33'b0100111100010000_1_0_xx_001_111_xxx_1_x_xx;
      patterns[9635] = 33'b0100111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9636] = 33'b0000011111010000_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9637] = 33'b0000111111010000_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9638] = 33'b0000111111010000_0_0_00_000_000_000_0_0_00;
      patterns[9639] = 33'b1000011100010011_0_1_00_001_011_111_0_x_00;
      patterns[9640] = 33'b1000111100010011_1_1_00_001_011_111_0_x_00;
      patterns[9641] = 33'b1000111100010011_0_0_00_000_000_000_0_0_00;
      patterns[9642] = 33'b1001011100010011_0_1_01_001_011_111_0_x_00;
      patterns[9643] = 33'b1001111100010011_1_1_01_001_011_111_0_x_00;
      patterns[9644] = 33'b1001111100010011_0_0_00_000_000_000_0_0_00;
      patterns[9645] = 33'b1010011100010011_0_1_10_001_011_111_0_x_00;
      patterns[9646] = 33'b1010111100010011_1_1_10_001_011_111_0_x_00;
      patterns[9647] = 33'b1010111100010011_0_0_00_000_000_000_0_0_00;
      patterns[9648] = 33'b1011011100010011_0_1_11_001_011_111_0_x_00;
      patterns[9649] = 33'b1011111100010011_1_1_11_001_011_111_0_x_00;
      patterns[9650] = 33'b1011111100010011_0_0_00_000_000_000_0_0_00;
      patterns[9651] = 33'b0101011100010000_0_1_xx_001_xxx_111_0_1_01;
      patterns[9652] = 33'b0101111100010000_1_1_xx_001_xxx_111_0_1_01;
      patterns[9653] = 33'b0101111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9654] = 33'b0100011100010000_0_0_xx_001_111_xxx_1_x_xx;
      patterns[9655] = 33'b0100111100010000_1_0_xx_001_111_xxx_1_x_xx;
      patterns[9656] = 33'b0100111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9657] = 33'b0000011100110100_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9658] = 33'b0000111100110100_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9659] = 33'b0000111100110100_0_0_00_000_000_000_0_0_00;
      patterns[9660] = 33'b1000011100010100_0_1_00_001_100_111_0_x_00;
      patterns[9661] = 33'b1000111100010100_1_1_00_001_100_111_0_x_00;
      patterns[9662] = 33'b1000111100010100_0_0_00_000_000_000_0_0_00;
      patterns[9663] = 33'b1001011100010100_0_1_01_001_100_111_0_x_00;
      patterns[9664] = 33'b1001111100010100_1_1_01_001_100_111_0_x_00;
      patterns[9665] = 33'b1001111100010100_0_0_00_000_000_000_0_0_00;
      patterns[9666] = 33'b1010011100010100_0_1_10_001_100_111_0_x_00;
      patterns[9667] = 33'b1010111100010100_1_1_10_001_100_111_0_x_00;
      patterns[9668] = 33'b1010111100010100_0_0_00_000_000_000_0_0_00;
      patterns[9669] = 33'b1011011100010100_0_1_11_001_100_111_0_x_00;
      patterns[9670] = 33'b1011111100010100_1_1_11_001_100_111_0_x_00;
      patterns[9671] = 33'b1011111100010100_0_0_00_000_000_000_0_0_00;
      patterns[9672] = 33'b0101011100010000_0_1_xx_001_xxx_111_0_1_01;
      patterns[9673] = 33'b0101111100010000_1_1_xx_001_xxx_111_0_1_01;
      patterns[9674] = 33'b0101111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9675] = 33'b0100011100010000_0_0_xx_001_111_xxx_1_x_xx;
      patterns[9676] = 33'b0100111100010000_1_0_xx_001_111_xxx_1_x_xx;
      patterns[9677] = 33'b0100111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9678] = 33'b0000011110001001_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9679] = 33'b0000111110001001_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9680] = 33'b0000111110001001_0_0_00_000_000_000_0_0_00;
      patterns[9681] = 33'b1000011100010101_0_1_00_001_101_111_0_x_00;
      patterns[9682] = 33'b1000111100010101_1_1_00_001_101_111_0_x_00;
      patterns[9683] = 33'b1000111100010101_0_0_00_000_000_000_0_0_00;
      patterns[9684] = 33'b1001011100010101_0_1_01_001_101_111_0_x_00;
      patterns[9685] = 33'b1001111100010101_1_1_01_001_101_111_0_x_00;
      patterns[9686] = 33'b1001111100010101_0_0_00_000_000_000_0_0_00;
      patterns[9687] = 33'b1010011100010101_0_1_10_001_101_111_0_x_00;
      patterns[9688] = 33'b1010111100010101_1_1_10_001_101_111_0_x_00;
      patterns[9689] = 33'b1010111100010101_0_0_00_000_000_000_0_0_00;
      patterns[9690] = 33'b1011011100010101_0_1_11_001_101_111_0_x_00;
      patterns[9691] = 33'b1011111100010101_1_1_11_001_101_111_0_x_00;
      patterns[9692] = 33'b1011111100010101_0_0_00_000_000_000_0_0_00;
      patterns[9693] = 33'b0101011100010000_0_1_xx_001_xxx_111_0_1_01;
      patterns[9694] = 33'b0101111100010000_1_1_xx_001_xxx_111_0_1_01;
      patterns[9695] = 33'b0101111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9696] = 33'b0100011100010000_0_0_xx_001_111_xxx_1_x_xx;
      patterns[9697] = 33'b0100111100010000_1_0_xx_001_111_xxx_1_x_xx;
      patterns[9698] = 33'b0100111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9699] = 33'b0000011110000111_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9700] = 33'b0000111110000111_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9701] = 33'b0000111110000111_0_0_00_000_000_000_0_0_00;
      patterns[9702] = 33'b1000011100010110_0_1_00_001_110_111_0_x_00;
      patterns[9703] = 33'b1000111100010110_1_1_00_001_110_111_0_x_00;
      patterns[9704] = 33'b1000111100010110_0_0_00_000_000_000_0_0_00;
      patterns[9705] = 33'b1001011100010110_0_1_01_001_110_111_0_x_00;
      patterns[9706] = 33'b1001111100010110_1_1_01_001_110_111_0_x_00;
      patterns[9707] = 33'b1001111100010110_0_0_00_000_000_000_0_0_00;
      patterns[9708] = 33'b1010011100010110_0_1_10_001_110_111_0_x_00;
      patterns[9709] = 33'b1010111100010110_1_1_10_001_110_111_0_x_00;
      patterns[9710] = 33'b1010111100010110_0_0_00_000_000_000_0_0_00;
      patterns[9711] = 33'b1011011100010110_0_1_11_001_110_111_0_x_00;
      patterns[9712] = 33'b1011111100010110_1_1_11_001_110_111_0_x_00;
      patterns[9713] = 33'b1011111100010110_0_0_00_000_000_000_0_0_00;
      patterns[9714] = 33'b0101011100010000_0_1_xx_001_xxx_111_0_1_01;
      patterns[9715] = 33'b0101111100010000_1_1_xx_001_xxx_111_0_1_01;
      patterns[9716] = 33'b0101111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9717] = 33'b0100011100010000_0_0_xx_001_111_xxx_1_x_xx;
      patterns[9718] = 33'b0100111100010000_1_0_xx_001_111_xxx_1_x_xx;
      patterns[9719] = 33'b0100111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9720] = 33'b0000011100101100_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9721] = 33'b0000111100101100_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9722] = 33'b0000111100101100_0_0_00_000_000_000_0_0_00;
      patterns[9723] = 33'b1000011100010111_0_1_00_001_111_111_0_x_00;
      patterns[9724] = 33'b1000111100010111_1_1_00_001_111_111_0_x_00;
      patterns[9725] = 33'b1000111100010111_0_0_00_000_000_000_0_0_00;
      patterns[9726] = 33'b1001011100010111_0_1_01_001_111_111_0_x_00;
      patterns[9727] = 33'b1001111100010111_1_1_01_001_111_111_0_x_00;
      patterns[9728] = 33'b1001111100010111_0_0_00_000_000_000_0_0_00;
      patterns[9729] = 33'b1010011100010111_0_1_10_001_111_111_0_x_00;
      patterns[9730] = 33'b1010111100010111_1_1_10_001_111_111_0_x_00;
      patterns[9731] = 33'b1010111100010111_0_0_00_000_000_000_0_0_00;
      patterns[9732] = 33'b1011011100010111_0_1_11_001_111_111_0_x_00;
      patterns[9733] = 33'b1011111100010111_1_1_11_001_111_111_0_x_00;
      patterns[9734] = 33'b1011111100010111_0_0_00_000_000_000_0_0_00;
      patterns[9735] = 33'b0101011100010000_0_1_xx_001_xxx_111_0_1_01;
      patterns[9736] = 33'b0101111100010000_1_1_xx_001_xxx_111_0_1_01;
      patterns[9737] = 33'b0101111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9738] = 33'b0100011100010000_0_0_xx_001_111_xxx_1_x_xx;
      patterns[9739] = 33'b0100111100010000_1_0_xx_001_111_xxx_1_x_xx;
      patterns[9740] = 33'b0100111100010000_0_0_00_000_000_000_0_0_00;
      patterns[9741] = 33'b0000011110001001_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9742] = 33'b0000111110001001_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9743] = 33'b0000111110001001_0_0_00_000_000_000_0_0_00;
      patterns[9744] = 33'b1000011100100000_0_1_00_010_000_111_0_x_00;
      patterns[9745] = 33'b1000111100100000_1_1_00_010_000_111_0_x_00;
      patterns[9746] = 33'b1000111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9747] = 33'b1001011100100000_0_1_01_010_000_111_0_x_00;
      patterns[9748] = 33'b1001111100100000_1_1_01_010_000_111_0_x_00;
      patterns[9749] = 33'b1001111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9750] = 33'b1010011100100000_0_1_10_010_000_111_0_x_00;
      patterns[9751] = 33'b1010111100100000_1_1_10_010_000_111_0_x_00;
      patterns[9752] = 33'b1010111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9753] = 33'b1011011100100000_0_1_11_010_000_111_0_x_00;
      patterns[9754] = 33'b1011111100100000_1_1_11_010_000_111_0_x_00;
      patterns[9755] = 33'b1011111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9756] = 33'b0101011100100000_0_1_xx_010_xxx_111_0_1_01;
      patterns[9757] = 33'b0101111100100000_1_1_xx_010_xxx_111_0_1_01;
      patterns[9758] = 33'b0101111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9759] = 33'b0100011100100000_0_0_xx_010_111_xxx_1_x_xx;
      patterns[9760] = 33'b0100111100100000_1_0_xx_010_111_xxx_1_x_xx;
      patterns[9761] = 33'b0100111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9762] = 33'b0000011111111100_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9763] = 33'b0000111111111100_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9764] = 33'b0000111111111100_0_0_00_000_000_000_0_0_00;
      patterns[9765] = 33'b1000011100100001_0_1_00_010_001_111_0_x_00;
      patterns[9766] = 33'b1000111100100001_1_1_00_010_001_111_0_x_00;
      patterns[9767] = 33'b1000111100100001_0_0_00_000_000_000_0_0_00;
      patterns[9768] = 33'b1001011100100001_0_1_01_010_001_111_0_x_00;
      patterns[9769] = 33'b1001111100100001_1_1_01_010_001_111_0_x_00;
      patterns[9770] = 33'b1001111100100001_0_0_00_000_000_000_0_0_00;
      patterns[9771] = 33'b1010011100100001_0_1_10_010_001_111_0_x_00;
      patterns[9772] = 33'b1010111100100001_1_1_10_010_001_111_0_x_00;
      patterns[9773] = 33'b1010111100100001_0_0_00_000_000_000_0_0_00;
      patterns[9774] = 33'b1011011100100001_0_1_11_010_001_111_0_x_00;
      patterns[9775] = 33'b1011111100100001_1_1_11_010_001_111_0_x_00;
      patterns[9776] = 33'b1011111100100001_0_0_00_000_000_000_0_0_00;
      patterns[9777] = 33'b0101011100100000_0_1_xx_010_xxx_111_0_1_01;
      patterns[9778] = 33'b0101111100100000_1_1_xx_010_xxx_111_0_1_01;
      patterns[9779] = 33'b0101111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9780] = 33'b0100011100100000_0_0_xx_010_111_xxx_1_x_xx;
      patterns[9781] = 33'b0100111100100000_1_0_xx_010_111_xxx_1_x_xx;
      patterns[9782] = 33'b0100111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9783] = 33'b0000011100111111_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9784] = 33'b0000111100111111_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9785] = 33'b0000111100111111_0_0_00_000_000_000_0_0_00;
      patterns[9786] = 33'b1000011100100010_0_1_00_010_010_111_0_x_00;
      patterns[9787] = 33'b1000111100100010_1_1_00_010_010_111_0_x_00;
      patterns[9788] = 33'b1000111100100010_0_0_00_000_000_000_0_0_00;
      patterns[9789] = 33'b1001011100100010_0_1_01_010_010_111_0_x_00;
      patterns[9790] = 33'b1001111100100010_1_1_01_010_010_111_0_x_00;
      patterns[9791] = 33'b1001111100100010_0_0_00_000_000_000_0_0_00;
      patterns[9792] = 33'b1010011100100010_0_1_10_010_010_111_0_x_00;
      patterns[9793] = 33'b1010111100100010_1_1_10_010_010_111_0_x_00;
      patterns[9794] = 33'b1010111100100010_0_0_00_000_000_000_0_0_00;
      patterns[9795] = 33'b1011011100100010_0_1_11_010_010_111_0_x_00;
      patterns[9796] = 33'b1011111100100010_1_1_11_010_010_111_0_x_00;
      patterns[9797] = 33'b1011111100100010_0_0_00_000_000_000_0_0_00;
      patterns[9798] = 33'b0101011100100000_0_1_xx_010_xxx_111_0_1_01;
      patterns[9799] = 33'b0101111100100000_1_1_xx_010_xxx_111_0_1_01;
      patterns[9800] = 33'b0101111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9801] = 33'b0100011100100000_0_0_xx_010_111_xxx_1_x_xx;
      patterns[9802] = 33'b0100111100100000_1_0_xx_010_111_xxx_1_x_xx;
      patterns[9803] = 33'b0100111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9804] = 33'b0000011111100000_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9805] = 33'b0000111111100000_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9806] = 33'b0000111111100000_0_0_00_000_000_000_0_0_00;
      patterns[9807] = 33'b1000011100100011_0_1_00_010_011_111_0_x_00;
      patterns[9808] = 33'b1000111100100011_1_1_00_010_011_111_0_x_00;
      patterns[9809] = 33'b1000111100100011_0_0_00_000_000_000_0_0_00;
      patterns[9810] = 33'b1001011100100011_0_1_01_010_011_111_0_x_00;
      patterns[9811] = 33'b1001111100100011_1_1_01_010_011_111_0_x_00;
      patterns[9812] = 33'b1001111100100011_0_0_00_000_000_000_0_0_00;
      patterns[9813] = 33'b1010011100100011_0_1_10_010_011_111_0_x_00;
      patterns[9814] = 33'b1010111100100011_1_1_10_010_011_111_0_x_00;
      patterns[9815] = 33'b1010111100100011_0_0_00_000_000_000_0_0_00;
      patterns[9816] = 33'b1011011100100011_0_1_11_010_011_111_0_x_00;
      patterns[9817] = 33'b1011111100100011_1_1_11_010_011_111_0_x_00;
      patterns[9818] = 33'b1011111100100011_0_0_00_000_000_000_0_0_00;
      patterns[9819] = 33'b0101011100100000_0_1_xx_010_xxx_111_0_1_01;
      patterns[9820] = 33'b0101111100100000_1_1_xx_010_xxx_111_0_1_01;
      patterns[9821] = 33'b0101111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9822] = 33'b0100011100100000_0_0_xx_010_111_xxx_1_x_xx;
      patterns[9823] = 33'b0100111100100000_1_0_xx_010_111_xxx_1_x_xx;
      patterns[9824] = 33'b0100111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9825] = 33'b0000011110010001_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9826] = 33'b0000111110010001_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9827] = 33'b0000111110010001_0_0_00_000_000_000_0_0_00;
      patterns[9828] = 33'b1000011100100100_0_1_00_010_100_111_0_x_00;
      patterns[9829] = 33'b1000111100100100_1_1_00_010_100_111_0_x_00;
      patterns[9830] = 33'b1000111100100100_0_0_00_000_000_000_0_0_00;
      patterns[9831] = 33'b1001011100100100_0_1_01_010_100_111_0_x_00;
      patterns[9832] = 33'b1001111100100100_1_1_01_010_100_111_0_x_00;
      patterns[9833] = 33'b1001111100100100_0_0_00_000_000_000_0_0_00;
      patterns[9834] = 33'b1010011100100100_0_1_10_010_100_111_0_x_00;
      patterns[9835] = 33'b1010111100100100_1_1_10_010_100_111_0_x_00;
      patterns[9836] = 33'b1010111100100100_0_0_00_000_000_000_0_0_00;
      patterns[9837] = 33'b1011011100100100_0_1_11_010_100_111_0_x_00;
      patterns[9838] = 33'b1011111100100100_1_1_11_010_100_111_0_x_00;
      patterns[9839] = 33'b1011111100100100_0_0_00_000_000_000_0_0_00;
      patterns[9840] = 33'b0101011100100000_0_1_xx_010_xxx_111_0_1_01;
      patterns[9841] = 33'b0101111100100000_1_1_xx_010_xxx_111_0_1_01;
      patterns[9842] = 33'b0101111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9843] = 33'b0100011100100000_0_0_xx_010_111_xxx_1_x_xx;
      patterns[9844] = 33'b0100111100100000_1_0_xx_010_111_xxx_1_x_xx;
      patterns[9845] = 33'b0100111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9846] = 33'b0000011111010001_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9847] = 33'b0000111111010001_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9848] = 33'b0000111111010001_0_0_00_000_000_000_0_0_00;
      patterns[9849] = 33'b1000011100100101_0_1_00_010_101_111_0_x_00;
      patterns[9850] = 33'b1000111100100101_1_1_00_010_101_111_0_x_00;
      patterns[9851] = 33'b1000111100100101_0_0_00_000_000_000_0_0_00;
      patterns[9852] = 33'b1001011100100101_0_1_01_010_101_111_0_x_00;
      patterns[9853] = 33'b1001111100100101_1_1_01_010_101_111_0_x_00;
      patterns[9854] = 33'b1001111100100101_0_0_00_000_000_000_0_0_00;
      patterns[9855] = 33'b1010011100100101_0_1_10_010_101_111_0_x_00;
      patterns[9856] = 33'b1010111100100101_1_1_10_010_101_111_0_x_00;
      patterns[9857] = 33'b1010111100100101_0_0_00_000_000_000_0_0_00;
      patterns[9858] = 33'b1011011100100101_0_1_11_010_101_111_0_x_00;
      patterns[9859] = 33'b1011111100100101_1_1_11_010_101_111_0_x_00;
      patterns[9860] = 33'b1011111100100101_0_0_00_000_000_000_0_0_00;
      patterns[9861] = 33'b0101011100100000_0_1_xx_010_xxx_111_0_1_01;
      patterns[9862] = 33'b0101111100100000_1_1_xx_010_xxx_111_0_1_01;
      patterns[9863] = 33'b0101111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9864] = 33'b0100011100100000_0_0_xx_010_111_xxx_1_x_xx;
      patterns[9865] = 33'b0100111100100000_1_0_xx_010_111_xxx_1_x_xx;
      patterns[9866] = 33'b0100111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9867] = 33'b0000011110100110_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9868] = 33'b0000111110100110_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9869] = 33'b0000111110100110_0_0_00_000_000_000_0_0_00;
      patterns[9870] = 33'b1000011100100110_0_1_00_010_110_111_0_x_00;
      patterns[9871] = 33'b1000111100100110_1_1_00_010_110_111_0_x_00;
      patterns[9872] = 33'b1000111100100110_0_0_00_000_000_000_0_0_00;
      patterns[9873] = 33'b1001011100100110_0_1_01_010_110_111_0_x_00;
      patterns[9874] = 33'b1001111100100110_1_1_01_010_110_111_0_x_00;
      patterns[9875] = 33'b1001111100100110_0_0_00_000_000_000_0_0_00;
      patterns[9876] = 33'b1010011100100110_0_1_10_010_110_111_0_x_00;
      patterns[9877] = 33'b1010111100100110_1_1_10_010_110_111_0_x_00;
      patterns[9878] = 33'b1010111100100110_0_0_00_000_000_000_0_0_00;
      patterns[9879] = 33'b1011011100100110_0_1_11_010_110_111_0_x_00;
      patterns[9880] = 33'b1011111100100110_1_1_11_010_110_111_0_x_00;
      patterns[9881] = 33'b1011111100100110_0_0_00_000_000_000_0_0_00;
      patterns[9882] = 33'b0101011100100000_0_1_xx_010_xxx_111_0_1_01;
      patterns[9883] = 33'b0101111100100000_1_1_xx_010_xxx_111_0_1_01;
      patterns[9884] = 33'b0101111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9885] = 33'b0100011100100000_0_0_xx_010_111_xxx_1_x_xx;
      patterns[9886] = 33'b0100111100100000_1_0_xx_010_111_xxx_1_x_xx;
      patterns[9887] = 33'b0100111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9888] = 33'b0000011110010111_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9889] = 33'b0000111110010111_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9890] = 33'b0000111110010111_0_0_00_000_000_000_0_0_00;
      patterns[9891] = 33'b1000011100100111_0_1_00_010_111_111_0_x_00;
      patterns[9892] = 33'b1000111100100111_1_1_00_010_111_111_0_x_00;
      patterns[9893] = 33'b1000111100100111_0_0_00_000_000_000_0_0_00;
      patterns[9894] = 33'b1001011100100111_0_1_01_010_111_111_0_x_00;
      patterns[9895] = 33'b1001111100100111_1_1_01_010_111_111_0_x_00;
      patterns[9896] = 33'b1001111100100111_0_0_00_000_000_000_0_0_00;
      patterns[9897] = 33'b1010011100100111_0_1_10_010_111_111_0_x_00;
      patterns[9898] = 33'b1010111100100111_1_1_10_010_111_111_0_x_00;
      patterns[9899] = 33'b1010111100100111_0_0_00_000_000_000_0_0_00;
      patterns[9900] = 33'b1011011100100111_0_1_11_010_111_111_0_x_00;
      patterns[9901] = 33'b1011111100100111_1_1_11_010_111_111_0_x_00;
      patterns[9902] = 33'b1011111100100111_0_0_00_000_000_000_0_0_00;
      patterns[9903] = 33'b0101011100100000_0_1_xx_010_xxx_111_0_1_01;
      patterns[9904] = 33'b0101111100100000_1_1_xx_010_xxx_111_0_1_01;
      patterns[9905] = 33'b0101111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9906] = 33'b0100011100100000_0_0_xx_010_111_xxx_1_x_xx;
      patterns[9907] = 33'b0100111100100000_1_0_xx_010_111_xxx_1_x_xx;
      patterns[9908] = 33'b0100111100100000_0_0_00_000_000_000_0_0_00;
      patterns[9909] = 33'b0000011101001100_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9910] = 33'b0000111101001100_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9911] = 33'b0000111101001100_0_0_00_000_000_000_0_0_00;
      patterns[9912] = 33'b1000011100110000_0_1_00_011_000_111_0_x_00;
      patterns[9913] = 33'b1000111100110000_1_1_00_011_000_111_0_x_00;
      patterns[9914] = 33'b1000111100110000_0_0_00_000_000_000_0_0_00;
      patterns[9915] = 33'b1001011100110000_0_1_01_011_000_111_0_x_00;
      patterns[9916] = 33'b1001111100110000_1_1_01_011_000_111_0_x_00;
      patterns[9917] = 33'b1001111100110000_0_0_00_000_000_000_0_0_00;
      patterns[9918] = 33'b1010011100110000_0_1_10_011_000_111_0_x_00;
      patterns[9919] = 33'b1010111100110000_1_1_10_011_000_111_0_x_00;
      patterns[9920] = 33'b1010111100110000_0_0_00_000_000_000_0_0_00;
      patterns[9921] = 33'b1011011100110000_0_1_11_011_000_111_0_x_00;
      patterns[9922] = 33'b1011111100110000_1_1_11_011_000_111_0_x_00;
      patterns[9923] = 33'b1011111100110000_0_0_00_000_000_000_0_0_00;
      patterns[9924] = 33'b0101011100110000_0_1_xx_011_xxx_111_0_1_01;
      patterns[9925] = 33'b0101111100110000_1_1_xx_011_xxx_111_0_1_01;
      patterns[9926] = 33'b0101111100110000_0_0_00_000_000_000_0_0_00;
      patterns[9927] = 33'b0100011100110000_0_0_xx_011_111_xxx_1_x_xx;
      patterns[9928] = 33'b0100111100110000_1_0_xx_011_111_xxx_1_x_xx;
      patterns[9929] = 33'b0100111100110000_0_0_00_000_000_000_0_0_00;
      patterns[9930] = 33'b0000011110010010_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9931] = 33'b0000111110010010_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9932] = 33'b0000111110010010_0_0_00_000_000_000_0_0_00;
      patterns[9933] = 33'b1000011100110001_0_1_00_011_001_111_0_x_00;
      patterns[9934] = 33'b1000111100110001_1_1_00_011_001_111_0_x_00;
      patterns[9935] = 33'b1000111100110001_0_0_00_000_000_000_0_0_00;
      patterns[9936] = 33'b1001011100110001_0_1_01_011_001_111_0_x_00;
      patterns[9937] = 33'b1001111100110001_1_1_01_011_001_111_0_x_00;
      patterns[9938] = 33'b1001111100110001_0_0_00_000_000_000_0_0_00;
      patterns[9939] = 33'b1010011100110001_0_1_10_011_001_111_0_x_00;
      patterns[9940] = 33'b1010111100110001_1_1_10_011_001_111_0_x_00;
      patterns[9941] = 33'b1010111100110001_0_0_00_000_000_000_0_0_00;
      patterns[9942] = 33'b1011011100110001_0_1_11_011_001_111_0_x_00;
      patterns[9943] = 33'b1011111100110001_1_1_11_011_001_111_0_x_00;
      patterns[9944] = 33'b1011111100110001_0_0_00_000_000_000_0_0_00;
      patterns[9945] = 33'b0101011100110000_0_1_xx_011_xxx_111_0_1_01;
      patterns[9946] = 33'b0101111100110000_1_1_xx_011_xxx_111_0_1_01;
      patterns[9947] = 33'b0101111100110000_0_0_00_000_000_000_0_0_00;
      patterns[9948] = 33'b0100011100110000_0_0_xx_011_111_xxx_1_x_xx;
      patterns[9949] = 33'b0100111100110000_1_0_xx_011_111_xxx_1_x_xx;
      patterns[9950] = 33'b0100111100110000_0_0_00_000_000_000_0_0_00;
      patterns[9951] = 33'b0000011101111011_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9952] = 33'b0000111101111011_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9953] = 33'b0000111101111011_0_0_00_000_000_000_0_0_00;
      patterns[9954] = 33'b1000011100110010_0_1_00_011_010_111_0_x_00;
      patterns[9955] = 33'b1000111100110010_1_1_00_011_010_111_0_x_00;
      patterns[9956] = 33'b1000111100110010_0_0_00_000_000_000_0_0_00;
      patterns[9957] = 33'b1001011100110010_0_1_01_011_010_111_0_x_00;
      patterns[9958] = 33'b1001111100110010_1_1_01_011_010_111_0_x_00;
      patterns[9959] = 33'b1001111100110010_0_0_00_000_000_000_0_0_00;
      patterns[9960] = 33'b1010011100110010_0_1_10_011_010_111_0_x_00;
      patterns[9961] = 33'b1010111100110010_1_1_10_011_010_111_0_x_00;
      patterns[9962] = 33'b1010111100110010_0_0_00_000_000_000_0_0_00;
      patterns[9963] = 33'b1011011100110010_0_1_11_011_010_111_0_x_00;
      patterns[9964] = 33'b1011111100110010_1_1_11_011_010_111_0_x_00;
      patterns[9965] = 33'b1011111100110010_0_0_00_000_000_000_0_0_00;
      patterns[9966] = 33'b0101011100110000_0_1_xx_011_xxx_111_0_1_01;
      patterns[9967] = 33'b0101111100110000_1_1_xx_011_xxx_111_0_1_01;
      patterns[9968] = 33'b0101111100110000_0_0_00_000_000_000_0_0_00;
      patterns[9969] = 33'b0100011100110000_0_0_xx_011_111_xxx_1_x_xx;
      patterns[9970] = 33'b0100111100110000_1_0_xx_011_111_xxx_1_x_xx;
      patterns[9971] = 33'b0100111100110000_0_0_00_000_000_000_0_0_00;
      patterns[9972] = 33'b0000011101101000_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9973] = 33'b0000111101101000_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9974] = 33'b0000111101101000_0_0_00_000_000_000_0_0_00;
      patterns[9975] = 33'b1000011100110011_0_1_00_011_011_111_0_x_00;
      patterns[9976] = 33'b1000111100110011_1_1_00_011_011_111_0_x_00;
      patterns[9977] = 33'b1000111100110011_0_0_00_000_000_000_0_0_00;
      patterns[9978] = 33'b1001011100110011_0_1_01_011_011_111_0_x_00;
      patterns[9979] = 33'b1001111100110011_1_1_01_011_011_111_0_x_00;
      patterns[9980] = 33'b1001111100110011_0_0_00_000_000_000_0_0_00;
      patterns[9981] = 33'b1010011100110011_0_1_10_011_011_111_0_x_00;
      patterns[9982] = 33'b1010111100110011_1_1_10_011_011_111_0_x_00;
      patterns[9983] = 33'b1010111100110011_0_0_00_000_000_000_0_0_00;
      patterns[9984] = 33'b1011011100110011_0_1_11_011_011_111_0_x_00;
      patterns[9985] = 33'b1011111100110011_1_1_11_011_011_111_0_x_00;
      patterns[9986] = 33'b1011111100110011_0_0_00_000_000_000_0_0_00;
      patterns[9987] = 33'b0101011100110000_0_1_xx_011_xxx_111_0_1_01;
      patterns[9988] = 33'b0101111100110000_1_1_xx_011_xxx_111_0_1_01;
      patterns[9989] = 33'b0101111100110000_0_0_00_000_000_000_0_0_00;
      patterns[9990] = 33'b0100011100110000_0_0_xx_011_111_xxx_1_x_xx;
      patterns[9991] = 33'b0100111100110000_1_0_xx_011_111_xxx_1_x_xx;
      patterns[9992] = 33'b0100111100110000_0_0_00_000_000_000_0_0_00;
      patterns[9993] = 33'b0000011111111111_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[9994] = 33'b0000111111111111_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[9995] = 33'b0000111111111111_0_0_00_000_000_000_0_0_00;
      patterns[9996] = 33'b1000011100110100_0_1_00_011_100_111_0_x_00;
      patterns[9997] = 33'b1000111100110100_1_1_00_011_100_111_0_x_00;
      patterns[9998] = 33'b1000111100110100_0_0_00_000_000_000_0_0_00;
      patterns[9999] = 33'b1001011100110100_0_1_01_011_100_111_0_x_00;
      patterns[10000] = 33'b1001111100110100_1_1_01_011_100_111_0_x_00;
      patterns[10001] = 33'b1001111100110100_0_0_00_000_000_000_0_0_00;
      patterns[10002] = 33'b1010011100110100_0_1_10_011_100_111_0_x_00;
      patterns[10003] = 33'b1010111100110100_1_1_10_011_100_111_0_x_00;
      patterns[10004] = 33'b1010111100110100_0_0_00_000_000_000_0_0_00;
      patterns[10005] = 33'b1011011100110100_0_1_11_011_100_111_0_x_00;
      patterns[10006] = 33'b1011111100110100_1_1_11_011_100_111_0_x_00;
      patterns[10007] = 33'b1011111100110100_0_0_00_000_000_000_0_0_00;
      patterns[10008] = 33'b0101011100110000_0_1_xx_011_xxx_111_0_1_01;
      patterns[10009] = 33'b0101111100110000_1_1_xx_011_xxx_111_0_1_01;
      patterns[10010] = 33'b0101111100110000_0_0_00_000_000_000_0_0_00;
      patterns[10011] = 33'b0100011100110000_0_0_xx_011_111_xxx_1_x_xx;
      patterns[10012] = 33'b0100111100110000_1_0_xx_011_111_xxx_1_x_xx;
      patterns[10013] = 33'b0100111100110000_0_0_00_000_000_000_0_0_00;
      patterns[10014] = 33'b0000011110011010_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10015] = 33'b0000111110011010_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10016] = 33'b0000111110011010_0_0_00_000_000_000_0_0_00;
      patterns[10017] = 33'b1000011100110101_0_1_00_011_101_111_0_x_00;
      patterns[10018] = 33'b1000111100110101_1_1_00_011_101_111_0_x_00;
      patterns[10019] = 33'b1000111100110101_0_0_00_000_000_000_0_0_00;
      patterns[10020] = 33'b1001011100110101_0_1_01_011_101_111_0_x_00;
      patterns[10021] = 33'b1001111100110101_1_1_01_011_101_111_0_x_00;
      patterns[10022] = 33'b1001111100110101_0_0_00_000_000_000_0_0_00;
      patterns[10023] = 33'b1010011100110101_0_1_10_011_101_111_0_x_00;
      patterns[10024] = 33'b1010111100110101_1_1_10_011_101_111_0_x_00;
      patterns[10025] = 33'b1010111100110101_0_0_00_000_000_000_0_0_00;
      patterns[10026] = 33'b1011011100110101_0_1_11_011_101_111_0_x_00;
      patterns[10027] = 33'b1011111100110101_1_1_11_011_101_111_0_x_00;
      patterns[10028] = 33'b1011111100110101_0_0_00_000_000_000_0_0_00;
      patterns[10029] = 33'b0101011100110000_0_1_xx_011_xxx_111_0_1_01;
      patterns[10030] = 33'b0101111100110000_1_1_xx_011_xxx_111_0_1_01;
      patterns[10031] = 33'b0101111100110000_0_0_00_000_000_000_0_0_00;
      patterns[10032] = 33'b0100011100110000_0_0_xx_011_111_xxx_1_x_xx;
      patterns[10033] = 33'b0100111100110000_1_0_xx_011_111_xxx_1_x_xx;
      patterns[10034] = 33'b0100111100110000_0_0_00_000_000_000_0_0_00;
      patterns[10035] = 33'b0000011101111001_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10036] = 33'b0000111101111001_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10037] = 33'b0000111101111001_0_0_00_000_000_000_0_0_00;
      patterns[10038] = 33'b1000011100110110_0_1_00_011_110_111_0_x_00;
      patterns[10039] = 33'b1000111100110110_1_1_00_011_110_111_0_x_00;
      patterns[10040] = 33'b1000111100110110_0_0_00_000_000_000_0_0_00;
      patterns[10041] = 33'b1001011100110110_0_1_01_011_110_111_0_x_00;
      patterns[10042] = 33'b1001111100110110_1_1_01_011_110_111_0_x_00;
      patterns[10043] = 33'b1001111100110110_0_0_00_000_000_000_0_0_00;
      patterns[10044] = 33'b1010011100110110_0_1_10_011_110_111_0_x_00;
      patterns[10045] = 33'b1010111100110110_1_1_10_011_110_111_0_x_00;
      patterns[10046] = 33'b1010111100110110_0_0_00_000_000_000_0_0_00;
      patterns[10047] = 33'b1011011100110110_0_1_11_011_110_111_0_x_00;
      patterns[10048] = 33'b1011111100110110_1_1_11_011_110_111_0_x_00;
      patterns[10049] = 33'b1011111100110110_0_0_00_000_000_000_0_0_00;
      patterns[10050] = 33'b0101011100110000_0_1_xx_011_xxx_111_0_1_01;
      patterns[10051] = 33'b0101111100110000_1_1_xx_011_xxx_111_0_1_01;
      patterns[10052] = 33'b0101111100110000_0_0_00_000_000_000_0_0_00;
      patterns[10053] = 33'b0100011100110000_0_0_xx_011_111_xxx_1_x_xx;
      patterns[10054] = 33'b0100111100110000_1_0_xx_011_111_xxx_1_x_xx;
      patterns[10055] = 33'b0100111100110000_0_0_00_000_000_000_0_0_00;
      patterns[10056] = 33'b0000011110101111_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10057] = 33'b0000111110101111_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10058] = 33'b0000111110101111_0_0_00_000_000_000_0_0_00;
      patterns[10059] = 33'b1000011100110111_0_1_00_011_111_111_0_x_00;
      patterns[10060] = 33'b1000111100110111_1_1_00_011_111_111_0_x_00;
      patterns[10061] = 33'b1000111100110111_0_0_00_000_000_000_0_0_00;
      patterns[10062] = 33'b1001011100110111_0_1_01_011_111_111_0_x_00;
      patterns[10063] = 33'b1001111100110111_1_1_01_011_111_111_0_x_00;
      patterns[10064] = 33'b1001111100110111_0_0_00_000_000_000_0_0_00;
      patterns[10065] = 33'b1010011100110111_0_1_10_011_111_111_0_x_00;
      patterns[10066] = 33'b1010111100110111_1_1_10_011_111_111_0_x_00;
      patterns[10067] = 33'b1010111100110111_0_0_00_000_000_000_0_0_00;
      patterns[10068] = 33'b1011011100110111_0_1_11_011_111_111_0_x_00;
      patterns[10069] = 33'b1011111100110111_1_1_11_011_111_111_0_x_00;
      patterns[10070] = 33'b1011111100110111_0_0_00_000_000_000_0_0_00;
      patterns[10071] = 33'b0101011100110000_0_1_xx_011_xxx_111_0_1_01;
      patterns[10072] = 33'b0101111100110000_1_1_xx_011_xxx_111_0_1_01;
      patterns[10073] = 33'b0101111100110000_0_0_00_000_000_000_0_0_00;
      patterns[10074] = 33'b0100011100110000_0_0_xx_011_111_xxx_1_x_xx;
      patterns[10075] = 33'b0100111100110000_1_0_xx_011_111_xxx_1_x_xx;
      patterns[10076] = 33'b0100111100110000_0_0_00_000_000_000_0_0_00;
      patterns[10077] = 33'b0000011111110100_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10078] = 33'b0000111111110100_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10079] = 33'b0000111111110100_0_0_00_000_000_000_0_0_00;
      patterns[10080] = 33'b1000011101000000_0_1_00_100_000_111_0_x_00;
      patterns[10081] = 33'b1000111101000000_1_1_00_100_000_111_0_x_00;
      patterns[10082] = 33'b1000111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10083] = 33'b1001011101000000_0_1_01_100_000_111_0_x_00;
      patterns[10084] = 33'b1001111101000000_1_1_01_100_000_111_0_x_00;
      patterns[10085] = 33'b1001111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10086] = 33'b1010011101000000_0_1_10_100_000_111_0_x_00;
      patterns[10087] = 33'b1010111101000000_1_1_10_100_000_111_0_x_00;
      patterns[10088] = 33'b1010111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10089] = 33'b1011011101000000_0_1_11_100_000_111_0_x_00;
      patterns[10090] = 33'b1011111101000000_1_1_11_100_000_111_0_x_00;
      patterns[10091] = 33'b1011111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10092] = 33'b0101011101000000_0_1_xx_100_xxx_111_0_1_01;
      patterns[10093] = 33'b0101111101000000_1_1_xx_100_xxx_111_0_1_01;
      patterns[10094] = 33'b0101111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10095] = 33'b0100011101000000_0_0_xx_100_111_xxx_1_x_xx;
      patterns[10096] = 33'b0100111101000000_1_0_xx_100_111_xxx_1_x_xx;
      patterns[10097] = 33'b0100111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10098] = 33'b0000011110101111_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10099] = 33'b0000111110101111_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10100] = 33'b0000111110101111_0_0_00_000_000_000_0_0_00;
      patterns[10101] = 33'b1000011101000001_0_1_00_100_001_111_0_x_00;
      patterns[10102] = 33'b1000111101000001_1_1_00_100_001_111_0_x_00;
      patterns[10103] = 33'b1000111101000001_0_0_00_000_000_000_0_0_00;
      patterns[10104] = 33'b1001011101000001_0_1_01_100_001_111_0_x_00;
      patterns[10105] = 33'b1001111101000001_1_1_01_100_001_111_0_x_00;
      patterns[10106] = 33'b1001111101000001_0_0_00_000_000_000_0_0_00;
      patterns[10107] = 33'b1010011101000001_0_1_10_100_001_111_0_x_00;
      patterns[10108] = 33'b1010111101000001_1_1_10_100_001_111_0_x_00;
      patterns[10109] = 33'b1010111101000001_0_0_00_000_000_000_0_0_00;
      patterns[10110] = 33'b1011011101000001_0_1_11_100_001_111_0_x_00;
      patterns[10111] = 33'b1011111101000001_1_1_11_100_001_111_0_x_00;
      patterns[10112] = 33'b1011111101000001_0_0_00_000_000_000_0_0_00;
      patterns[10113] = 33'b0101011101000000_0_1_xx_100_xxx_111_0_1_01;
      patterns[10114] = 33'b0101111101000000_1_1_xx_100_xxx_111_0_1_01;
      patterns[10115] = 33'b0101111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10116] = 33'b0100011101000000_0_0_xx_100_111_xxx_1_x_xx;
      patterns[10117] = 33'b0100111101000000_1_0_xx_100_111_xxx_1_x_xx;
      patterns[10118] = 33'b0100111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10119] = 33'b0000011101010100_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10120] = 33'b0000111101010100_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10121] = 33'b0000111101010100_0_0_00_000_000_000_0_0_00;
      patterns[10122] = 33'b1000011101000010_0_1_00_100_010_111_0_x_00;
      patterns[10123] = 33'b1000111101000010_1_1_00_100_010_111_0_x_00;
      patterns[10124] = 33'b1000111101000010_0_0_00_000_000_000_0_0_00;
      patterns[10125] = 33'b1001011101000010_0_1_01_100_010_111_0_x_00;
      patterns[10126] = 33'b1001111101000010_1_1_01_100_010_111_0_x_00;
      patterns[10127] = 33'b1001111101000010_0_0_00_000_000_000_0_0_00;
      patterns[10128] = 33'b1010011101000010_0_1_10_100_010_111_0_x_00;
      patterns[10129] = 33'b1010111101000010_1_1_10_100_010_111_0_x_00;
      patterns[10130] = 33'b1010111101000010_0_0_00_000_000_000_0_0_00;
      patterns[10131] = 33'b1011011101000010_0_1_11_100_010_111_0_x_00;
      patterns[10132] = 33'b1011111101000010_1_1_11_100_010_111_0_x_00;
      patterns[10133] = 33'b1011111101000010_0_0_00_000_000_000_0_0_00;
      patterns[10134] = 33'b0101011101000000_0_1_xx_100_xxx_111_0_1_01;
      patterns[10135] = 33'b0101111101000000_1_1_xx_100_xxx_111_0_1_01;
      patterns[10136] = 33'b0101111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10137] = 33'b0100011101000000_0_0_xx_100_111_xxx_1_x_xx;
      patterns[10138] = 33'b0100111101000000_1_0_xx_100_111_xxx_1_x_xx;
      patterns[10139] = 33'b0100111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10140] = 33'b0000011111100100_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10141] = 33'b0000111111100100_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10142] = 33'b0000111111100100_0_0_00_000_000_000_0_0_00;
      patterns[10143] = 33'b1000011101000011_0_1_00_100_011_111_0_x_00;
      patterns[10144] = 33'b1000111101000011_1_1_00_100_011_111_0_x_00;
      patterns[10145] = 33'b1000111101000011_0_0_00_000_000_000_0_0_00;
      patterns[10146] = 33'b1001011101000011_0_1_01_100_011_111_0_x_00;
      patterns[10147] = 33'b1001111101000011_1_1_01_100_011_111_0_x_00;
      patterns[10148] = 33'b1001111101000011_0_0_00_000_000_000_0_0_00;
      patterns[10149] = 33'b1010011101000011_0_1_10_100_011_111_0_x_00;
      patterns[10150] = 33'b1010111101000011_1_1_10_100_011_111_0_x_00;
      patterns[10151] = 33'b1010111101000011_0_0_00_000_000_000_0_0_00;
      patterns[10152] = 33'b1011011101000011_0_1_11_100_011_111_0_x_00;
      patterns[10153] = 33'b1011111101000011_1_1_11_100_011_111_0_x_00;
      patterns[10154] = 33'b1011111101000011_0_0_00_000_000_000_0_0_00;
      patterns[10155] = 33'b0101011101000000_0_1_xx_100_xxx_111_0_1_01;
      patterns[10156] = 33'b0101111101000000_1_1_xx_100_xxx_111_0_1_01;
      patterns[10157] = 33'b0101111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10158] = 33'b0100011101000000_0_0_xx_100_111_xxx_1_x_xx;
      patterns[10159] = 33'b0100111101000000_1_0_xx_100_111_xxx_1_x_xx;
      patterns[10160] = 33'b0100111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10161] = 33'b0000011110110111_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10162] = 33'b0000111110110111_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10163] = 33'b0000111110110111_0_0_00_000_000_000_0_0_00;
      patterns[10164] = 33'b1000011101000100_0_1_00_100_100_111_0_x_00;
      patterns[10165] = 33'b1000111101000100_1_1_00_100_100_111_0_x_00;
      patterns[10166] = 33'b1000111101000100_0_0_00_000_000_000_0_0_00;
      patterns[10167] = 33'b1001011101000100_0_1_01_100_100_111_0_x_00;
      patterns[10168] = 33'b1001111101000100_1_1_01_100_100_111_0_x_00;
      patterns[10169] = 33'b1001111101000100_0_0_00_000_000_000_0_0_00;
      patterns[10170] = 33'b1010011101000100_0_1_10_100_100_111_0_x_00;
      patterns[10171] = 33'b1010111101000100_1_1_10_100_100_111_0_x_00;
      patterns[10172] = 33'b1010111101000100_0_0_00_000_000_000_0_0_00;
      patterns[10173] = 33'b1011011101000100_0_1_11_100_100_111_0_x_00;
      patterns[10174] = 33'b1011111101000100_1_1_11_100_100_111_0_x_00;
      patterns[10175] = 33'b1011111101000100_0_0_00_000_000_000_0_0_00;
      patterns[10176] = 33'b0101011101000000_0_1_xx_100_xxx_111_0_1_01;
      patterns[10177] = 33'b0101111101000000_1_1_xx_100_xxx_111_0_1_01;
      patterns[10178] = 33'b0101111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10179] = 33'b0100011101000000_0_0_xx_100_111_xxx_1_x_xx;
      patterns[10180] = 33'b0100111101000000_1_0_xx_100_111_xxx_1_x_xx;
      patterns[10181] = 33'b0100111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10182] = 33'b0000011111001000_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10183] = 33'b0000111111001000_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10184] = 33'b0000111111001000_0_0_00_000_000_000_0_0_00;
      patterns[10185] = 33'b1000011101000101_0_1_00_100_101_111_0_x_00;
      patterns[10186] = 33'b1000111101000101_1_1_00_100_101_111_0_x_00;
      patterns[10187] = 33'b1000111101000101_0_0_00_000_000_000_0_0_00;
      patterns[10188] = 33'b1001011101000101_0_1_01_100_101_111_0_x_00;
      patterns[10189] = 33'b1001111101000101_1_1_01_100_101_111_0_x_00;
      patterns[10190] = 33'b1001111101000101_0_0_00_000_000_000_0_0_00;
      patterns[10191] = 33'b1010011101000101_0_1_10_100_101_111_0_x_00;
      patterns[10192] = 33'b1010111101000101_1_1_10_100_101_111_0_x_00;
      patterns[10193] = 33'b1010111101000101_0_0_00_000_000_000_0_0_00;
      patterns[10194] = 33'b1011011101000101_0_1_11_100_101_111_0_x_00;
      patterns[10195] = 33'b1011111101000101_1_1_11_100_101_111_0_x_00;
      patterns[10196] = 33'b1011111101000101_0_0_00_000_000_000_0_0_00;
      patterns[10197] = 33'b0101011101000000_0_1_xx_100_xxx_111_0_1_01;
      patterns[10198] = 33'b0101111101000000_1_1_xx_100_xxx_111_0_1_01;
      patterns[10199] = 33'b0101111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10200] = 33'b0100011101000000_0_0_xx_100_111_xxx_1_x_xx;
      patterns[10201] = 33'b0100111101000000_1_0_xx_100_111_xxx_1_x_xx;
      patterns[10202] = 33'b0100111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10203] = 33'b0000011110001111_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10204] = 33'b0000111110001111_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10205] = 33'b0000111110001111_0_0_00_000_000_000_0_0_00;
      patterns[10206] = 33'b1000011101000110_0_1_00_100_110_111_0_x_00;
      patterns[10207] = 33'b1000111101000110_1_1_00_100_110_111_0_x_00;
      patterns[10208] = 33'b1000111101000110_0_0_00_000_000_000_0_0_00;
      patterns[10209] = 33'b1001011101000110_0_1_01_100_110_111_0_x_00;
      patterns[10210] = 33'b1001111101000110_1_1_01_100_110_111_0_x_00;
      patterns[10211] = 33'b1001111101000110_0_0_00_000_000_000_0_0_00;
      patterns[10212] = 33'b1010011101000110_0_1_10_100_110_111_0_x_00;
      patterns[10213] = 33'b1010111101000110_1_1_10_100_110_111_0_x_00;
      patterns[10214] = 33'b1010111101000110_0_0_00_000_000_000_0_0_00;
      patterns[10215] = 33'b1011011101000110_0_1_11_100_110_111_0_x_00;
      patterns[10216] = 33'b1011111101000110_1_1_11_100_110_111_0_x_00;
      patterns[10217] = 33'b1011111101000110_0_0_00_000_000_000_0_0_00;
      patterns[10218] = 33'b0101011101000000_0_1_xx_100_xxx_111_0_1_01;
      patterns[10219] = 33'b0101111101000000_1_1_xx_100_xxx_111_0_1_01;
      patterns[10220] = 33'b0101111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10221] = 33'b0100011101000000_0_0_xx_100_111_xxx_1_x_xx;
      patterns[10222] = 33'b0100111101000000_1_0_xx_100_111_xxx_1_x_xx;
      patterns[10223] = 33'b0100111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10224] = 33'b0000011101010010_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10225] = 33'b0000111101010010_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10226] = 33'b0000111101010010_0_0_00_000_000_000_0_0_00;
      patterns[10227] = 33'b1000011101000111_0_1_00_100_111_111_0_x_00;
      patterns[10228] = 33'b1000111101000111_1_1_00_100_111_111_0_x_00;
      patterns[10229] = 33'b1000111101000111_0_0_00_000_000_000_0_0_00;
      patterns[10230] = 33'b1001011101000111_0_1_01_100_111_111_0_x_00;
      patterns[10231] = 33'b1001111101000111_1_1_01_100_111_111_0_x_00;
      patterns[10232] = 33'b1001111101000111_0_0_00_000_000_000_0_0_00;
      patterns[10233] = 33'b1010011101000111_0_1_10_100_111_111_0_x_00;
      patterns[10234] = 33'b1010111101000111_1_1_10_100_111_111_0_x_00;
      patterns[10235] = 33'b1010111101000111_0_0_00_000_000_000_0_0_00;
      patterns[10236] = 33'b1011011101000111_0_1_11_100_111_111_0_x_00;
      patterns[10237] = 33'b1011111101000111_1_1_11_100_111_111_0_x_00;
      patterns[10238] = 33'b1011111101000111_0_0_00_000_000_000_0_0_00;
      patterns[10239] = 33'b0101011101000000_0_1_xx_100_xxx_111_0_1_01;
      patterns[10240] = 33'b0101111101000000_1_1_xx_100_xxx_111_0_1_01;
      patterns[10241] = 33'b0101111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10242] = 33'b0100011101000000_0_0_xx_100_111_xxx_1_x_xx;
      patterns[10243] = 33'b0100111101000000_1_0_xx_100_111_xxx_1_x_xx;
      patterns[10244] = 33'b0100111101000000_0_0_00_000_000_000_0_0_00;
      patterns[10245] = 33'b0000011111101010_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10246] = 33'b0000111111101010_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10247] = 33'b0000111111101010_0_0_00_000_000_000_0_0_00;
      patterns[10248] = 33'b1000011101010000_0_1_00_101_000_111_0_x_00;
      patterns[10249] = 33'b1000111101010000_1_1_00_101_000_111_0_x_00;
      patterns[10250] = 33'b1000111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10251] = 33'b1001011101010000_0_1_01_101_000_111_0_x_00;
      patterns[10252] = 33'b1001111101010000_1_1_01_101_000_111_0_x_00;
      patterns[10253] = 33'b1001111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10254] = 33'b1010011101010000_0_1_10_101_000_111_0_x_00;
      patterns[10255] = 33'b1010111101010000_1_1_10_101_000_111_0_x_00;
      patterns[10256] = 33'b1010111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10257] = 33'b1011011101010000_0_1_11_101_000_111_0_x_00;
      patterns[10258] = 33'b1011111101010000_1_1_11_101_000_111_0_x_00;
      patterns[10259] = 33'b1011111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10260] = 33'b0101011101010000_0_1_xx_101_xxx_111_0_1_01;
      patterns[10261] = 33'b0101111101010000_1_1_xx_101_xxx_111_0_1_01;
      patterns[10262] = 33'b0101111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10263] = 33'b0100011101010000_0_0_xx_101_111_xxx_1_x_xx;
      patterns[10264] = 33'b0100111101010000_1_0_xx_101_111_xxx_1_x_xx;
      patterns[10265] = 33'b0100111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10266] = 33'b0000011110011111_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10267] = 33'b0000111110011111_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10268] = 33'b0000111110011111_0_0_00_000_000_000_0_0_00;
      patterns[10269] = 33'b1000011101010001_0_1_00_101_001_111_0_x_00;
      patterns[10270] = 33'b1000111101010001_1_1_00_101_001_111_0_x_00;
      patterns[10271] = 33'b1000111101010001_0_0_00_000_000_000_0_0_00;
      patterns[10272] = 33'b1001011101010001_0_1_01_101_001_111_0_x_00;
      patterns[10273] = 33'b1001111101010001_1_1_01_101_001_111_0_x_00;
      patterns[10274] = 33'b1001111101010001_0_0_00_000_000_000_0_0_00;
      patterns[10275] = 33'b1010011101010001_0_1_10_101_001_111_0_x_00;
      patterns[10276] = 33'b1010111101010001_1_1_10_101_001_111_0_x_00;
      patterns[10277] = 33'b1010111101010001_0_0_00_000_000_000_0_0_00;
      patterns[10278] = 33'b1011011101010001_0_1_11_101_001_111_0_x_00;
      patterns[10279] = 33'b1011111101010001_1_1_11_101_001_111_0_x_00;
      patterns[10280] = 33'b1011111101010001_0_0_00_000_000_000_0_0_00;
      patterns[10281] = 33'b0101011101010000_0_1_xx_101_xxx_111_0_1_01;
      patterns[10282] = 33'b0101111101010000_1_1_xx_101_xxx_111_0_1_01;
      patterns[10283] = 33'b0101111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10284] = 33'b0100011101010000_0_0_xx_101_111_xxx_1_x_xx;
      patterns[10285] = 33'b0100111101010000_1_0_xx_101_111_xxx_1_x_xx;
      patterns[10286] = 33'b0100111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10287] = 33'b0000011100111000_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10288] = 33'b0000111100111000_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10289] = 33'b0000111100111000_0_0_00_000_000_000_0_0_00;
      patterns[10290] = 33'b1000011101010010_0_1_00_101_010_111_0_x_00;
      patterns[10291] = 33'b1000111101010010_1_1_00_101_010_111_0_x_00;
      patterns[10292] = 33'b1000111101010010_0_0_00_000_000_000_0_0_00;
      patterns[10293] = 33'b1001011101010010_0_1_01_101_010_111_0_x_00;
      patterns[10294] = 33'b1001111101010010_1_1_01_101_010_111_0_x_00;
      patterns[10295] = 33'b1001111101010010_0_0_00_000_000_000_0_0_00;
      patterns[10296] = 33'b1010011101010010_0_1_10_101_010_111_0_x_00;
      patterns[10297] = 33'b1010111101010010_1_1_10_101_010_111_0_x_00;
      patterns[10298] = 33'b1010111101010010_0_0_00_000_000_000_0_0_00;
      patterns[10299] = 33'b1011011101010010_0_1_11_101_010_111_0_x_00;
      patterns[10300] = 33'b1011111101010010_1_1_11_101_010_111_0_x_00;
      patterns[10301] = 33'b1011111101010010_0_0_00_000_000_000_0_0_00;
      patterns[10302] = 33'b0101011101010000_0_1_xx_101_xxx_111_0_1_01;
      patterns[10303] = 33'b0101111101010000_1_1_xx_101_xxx_111_0_1_01;
      patterns[10304] = 33'b0101111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10305] = 33'b0100011101010000_0_0_xx_101_111_xxx_1_x_xx;
      patterns[10306] = 33'b0100111101010000_1_0_xx_101_111_xxx_1_x_xx;
      patterns[10307] = 33'b0100111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10308] = 33'b0000011110110010_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10309] = 33'b0000111110110010_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10310] = 33'b0000111110110010_0_0_00_000_000_000_0_0_00;
      patterns[10311] = 33'b1000011101010011_0_1_00_101_011_111_0_x_00;
      patterns[10312] = 33'b1000111101010011_1_1_00_101_011_111_0_x_00;
      patterns[10313] = 33'b1000111101010011_0_0_00_000_000_000_0_0_00;
      patterns[10314] = 33'b1001011101010011_0_1_01_101_011_111_0_x_00;
      patterns[10315] = 33'b1001111101010011_1_1_01_101_011_111_0_x_00;
      patterns[10316] = 33'b1001111101010011_0_0_00_000_000_000_0_0_00;
      patterns[10317] = 33'b1010011101010011_0_1_10_101_011_111_0_x_00;
      patterns[10318] = 33'b1010111101010011_1_1_10_101_011_111_0_x_00;
      patterns[10319] = 33'b1010111101010011_0_0_00_000_000_000_0_0_00;
      patterns[10320] = 33'b1011011101010011_0_1_11_101_011_111_0_x_00;
      patterns[10321] = 33'b1011111101010011_1_1_11_101_011_111_0_x_00;
      patterns[10322] = 33'b1011111101010011_0_0_00_000_000_000_0_0_00;
      patterns[10323] = 33'b0101011101010000_0_1_xx_101_xxx_111_0_1_01;
      patterns[10324] = 33'b0101111101010000_1_1_xx_101_xxx_111_0_1_01;
      patterns[10325] = 33'b0101111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10326] = 33'b0100011101010000_0_0_xx_101_111_xxx_1_x_xx;
      patterns[10327] = 33'b0100111101010000_1_0_xx_101_111_xxx_1_x_xx;
      patterns[10328] = 33'b0100111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10329] = 33'b0000011111000111_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10330] = 33'b0000111111000111_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10331] = 33'b0000111111000111_0_0_00_000_000_000_0_0_00;
      patterns[10332] = 33'b1000011101010100_0_1_00_101_100_111_0_x_00;
      patterns[10333] = 33'b1000111101010100_1_1_00_101_100_111_0_x_00;
      patterns[10334] = 33'b1000111101010100_0_0_00_000_000_000_0_0_00;
      patterns[10335] = 33'b1001011101010100_0_1_01_101_100_111_0_x_00;
      patterns[10336] = 33'b1001111101010100_1_1_01_101_100_111_0_x_00;
      patterns[10337] = 33'b1001111101010100_0_0_00_000_000_000_0_0_00;
      patterns[10338] = 33'b1010011101010100_0_1_10_101_100_111_0_x_00;
      patterns[10339] = 33'b1010111101010100_1_1_10_101_100_111_0_x_00;
      patterns[10340] = 33'b1010111101010100_0_0_00_000_000_000_0_0_00;
      patterns[10341] = 33'b1011011101010100_0_1_11_101_100_111_0_x_00;
      patterns[10342] = 33'b1011111101010100_1_1_11_101_100_111_0_x_00;
      patterns[10343] = 33'b1011111101010100_0_0_00_000_000_000_0_0_00;
      patterns[10344] = 33'b0101011101010000_0_1_xx_101_xxx_111_0_1_01;
      patterns[10345] = 33'b0101111101010000_1_1_xx_101_xxx_111_0_1_01;
      patterns[10346] = 33'b0101111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10347] = 33'b0100011101010000_0_0_xx_101_111_xxx_1_x_xx;
      patterns[10348] = 33'b0100111101010000_1_0_xx_101_111_xxx_1_x_xx;
      patterns[10349] = 33'b0100111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10350] = 33'b0000011101000101_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10351] = 33'b0000111101000101_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10352] = 33'b0000111101000101_0_0_00_000_000_000_0_0_00;
      patterns[10353] = 33'b1000011101010101_0_1_00_101_101_111_0_x_00;
      patterns[10354] = 33'b1000111101010101_1_1_00_101_101_111_0_x_00;
      patterns[10355] = 33'b1000111101010101_0_0_00_000_000_000_0_0_00;
      patterns[10356] = 33'b1001011101010101_0_1_01_101_101_111_0_x_00;
      patterns[10357] = 33'b1001111101010101_1_1_01_101_101_111_0_x_00;
      patterns[10358] = 33'b1001111101010101_0_0_00_000_000_000_0_0_00;
      patterns[10359] = 33'b1010011101010101_0_1_10_101_101_111_0_x_00;
      patterns[10360] = 33'b1010111101010101_1_1_10_101_101_111_0_x_00;
      patterns[10361] = 33'b1010111101010101_0_0_00_000_000_000_0_0_00;
      patterns[10362] = 33'b1011011101010101_0_1_11_101_101_111_0_x_00;
      patterns[10363] = 33'b1011111101010101_1_1_11_101_101_111_0_x_00;
      patterns[10364] = 33'b1011111101010101_0_0_00_000_000_000_0_0_00;
      patterns[10365] = 33'b0101011101010000_0_1_xx_101_xxx_111_0_1_01;
      patterns[10366] = 33'b0101111101010000_1_1_xx_101_xxx_111_0_1_01;
      patterns[10367] = 33'b0101111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10368] = 33'b0100011101010000_0_0_xx_101_111_xxx_1_x_xx;
      patterns[10369] = 33'b0100111101010000_1_0_xx_101_111_xxx_1_x_xx;
      patterns[10370] = 33'b0100111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10371] = 33'b0000011111010010_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10372] = 33'b0000111111010010_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10373] = 33'b0000111111010010_0_0_00_000_000_000_0_0_00;
      patterns[10374] = 33'b1000011101010110_0_1_00_101_110_111_0_x_00;
      patterns[10375] = 33'b1000111101010110_1_1_00_101_110_111_0_x_00;
      patterns[10376] = 33'b1000111101010110_0_0_00_000_000_000_0_0_00;
      patterns[10377] = 33'b1001011101010110_0_1_01_101_110_111_0_x_00;
      patterns[10378] = 33'b1001111101010110_1_1_01_101_110_111_0_x_00;
      patterns[10379] = 33'b1001111101010110_0_0_00_000_000_000_0_0_00;
      patterns[10380] = 33'b1010011101010110_0_1_10_101_110_111_0_x_00;
      patterns[10381] = 33'b1010111101010110_1_1_10_101_110_111_0_x_00;
      patterns[10382] = 33'b1010111101010110_0_0_00_000_000_000_0_0_00;
      patterns[10383] = 33'b1011011101010110_0_1_11_101_110_111_0_x_00;
      patterns[10384] = 33'b1011111101010110_1_1_11_101_110_111_0_x_00;
      patterns[10385] = 33'b1011111101010110_0_0_00_000_000_000_0_0_00;
      patterns[10386] = 33'b0101011101010000_0_1_xx_101_xxx_111_0_1_01;
      patterns[10387] = 33'b0101111101010000_1_1_xx_101_xxx_111_0_1_01;
      patterns[10388] = 33'b0101111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10389] = 33'b0100011101010000_0_0_xx_101_111_xxx_1_x_xx;
      patterns[10390] = 33'b0100111101010000_1_0_xx_101_111_xxx_1_x_xx;
      patterns[10391] = 33'b0100111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10392] = 33'b0000011111011010_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10393] = 33'b0000111111011010_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10394] = 33'b0000111111011010_0_0_00_000_000_000_0_0_00;
      patterns[10395] = 33'b1000011101010111_0_1_00_101_111_111_0_x_00;
      patterns[10396] = 33'b1000111101010111_1_1_00_101_111_111_0_x_00;
      patterns[10397] = 33'b1000111101010111_0_0_00_000_000_000_0_0_00;
      patterns[10398] = 33'b1001011101010111_0_1_01_101_111_111_0_x_00;
      patterns[10399] = 33'b1001111101010111_1_1_01_101_111_111_0_x_00;
      patterns[10400] = 33'b1001111101010111_0_0_00_000_000_000_0_0_00;
      patterns[10401] = 33'b1010011101010111_0_1_10_101_111_111_0_x_00;
      patterns[10402] = 33'b1010111101010111_1_1_10_101_111_111_0_x_00;
      patterns[10403] = 33'b1010111101010111_0_0_00_000_000_000_0_0_00;
      patterns[10404] = 33'b1011011101010111_0_1_11_101_111_111_0_x_00;
      patterns[10405] = 33'b1011111101010111_1_1_11_101_111_111_0_x_00;
      patterns[10406] = 33'b1011111101010111_0_0_00_000_000_000_0_0_00;
      patterns[10407] = 33'b0101011101010000_0_1_xx_101_xxx_111_0_1_01;
      patterns[10408] = 33'b0101111101010000_1_1_xx_101_xxx_111_0_1_01;
      patterns[10409] = 33'b0101111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10410] = 33'b0100011101010000_0_0_xx_101_111_xxx_1_x_xx;
      patterns[10411] = 33'b0100111101010000_1_0_xx_101_111_xxx_1_x_xx;
      patterns[10412] = 33'b0100111101010000_0_0_00_000_000_000_0_0_00;
      patterns[10413] = 33'b0000011110110111_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10414] = 33'b0000111110110111_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10415] = 33'b0000111110110111_0_0_00_000_000_000_0_0_00;
      patterns[10416] = 33'b1000011101100000_0_1_00_110_000_111_0_x_00;
      patterns[10417] = 33'b1000111101100000_1_1_00_110_000_111_0_x_00;
      patterns[10418] = 33'b1000111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10419] = 33'b1001011101100000_0_1_01_110_000_111_0_x_00;
      patterns[10420] = 33'b1001111101100000_1_1_01_110_000_111_0_x_00;
      patterns[10421] = 33'b1001111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10422] = 33'b1010011101100000_0_1_10_110_000_111_0_x_00;
      patterns[10423] = 33'b1010111101100000_1_1_10_110_000_111_0_x_00;
      patterns[10424] = 33'b1010111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10425] = 33'b1011011101100000_0_1_11_110_000_111_0_x_00;
      patterns[10426] = 33'b1011111101100000_1_1_11_110_000_111_0_x_00;
      patterns[10427] = 33'b1011111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10428] = 33'b0101011101100000_0_1_xx_110_xxx_111_0_1_01;
      patterns[10429] = 33'b0101111101100000_1_1_xx_110_xxx_111_0_1_01;
      patterns[10430] = 33'b0101111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10431] = 33'b0100011101100000_0_0_xx_110_111_xxx_1_x_xx;
      patterns[10432] = 33'b0100111101100000_1_0_xx_110_111_xxx_1_x_xx;
      patterns[10433] = 33'b0100111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10434] = 33'b0000011111010100_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10435] = 33'b0000111111010100_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10436] = 33'b0000111111010100_0_0_00_000_000_000_0_0_00;
      patterns[10437] = 33'b1000011101100001_0_1_00_110_001_111_0_x_00;
      patterns[10438] = 33'b1000111101100001_1_1_00_110_001_111_0_x_00;
      patterns[10439] = 33'b1000111101100001_0_0_00_000_000_000_0_0_00;
      patterns[10440] = 33'b1001011101100001_0_1_01_110_001_111_0_x_00;
      patterns[10441] = 33'b1001111101100001_1_1_01_110_001_111_0_x_00;
      patterns[10442] = 33'b1001111101100001_0_0_00_000_000_000_0_0_00;
      patterns[10443] = 33'b1010011101100001_0_1_10_110_001_111_0_x_00;
      patterns[10444] = 33'b1010111101100001_1_1_10_110_001_111_0_x_00;
      patterns[10445] = 33'b1010111101100001_0_0_00_000_000_000_0_0_00;
      patterns[10446] = 33'b1011011101100001_0_1_11_110_001_111_0_x_00;
      patterns[10447] = 33'b1011111101100001_1_1_11_110_001_111_0_x_00;
      patterns[10448] = 33'b1011111101100001_0_0_00_000_000_000_0_0_00;
      patterns[10449] = 33'b0101011101100000_0_1_xx_110_xxx_111_0_1_01;
      patterns[10450] = 33'b0101111101100000_1_1_xx_110_xxx_111_0_1_01;
      patterns[10451] = 33'b0101111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10452] = 33'b0100011101100000_0_0_xx_110_111_xxx_1_x_xx;
      patterns[10453] = 33'b0100111101100000_1_0_xx_110_111_xxx_1_x_xx;
      patterns[10454] = 33'b0100111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10455] = 33'b0000011100010011_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10456] = 33'b0000111100010011_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10457] = 33'b0000111100010011_0_0_00_000_000_000_0_0_00;
      patterns[10458] = 33'b1000011101100010_0_1_00_110_010_111_0_x_00;
      patterns[10459] = 33'b1000111101100010_1_1_00_110_010_111_0_x_00;
      patterns[10460] = 33'b1000111101100010_0_0_00_000_000_000_0_0_00;
      patterns[10461] = 33'b1001011101100010_0_1_01_110_010_111_0_x_00;
      patterns[10462] = 33'b1001111101100010_1_1_01_110_010_111_0_x_00;
      patterns[10463] = 33'b1001111101100010_0_0_00_000_000_000_0_0_00;
      patterns[10464] = 33'b1010011101100010_0_1_10_110_010_111_0_x_00;
      patterns[10465] = 33'b1010111101100010_1_1_10_110_010_111_0_x_00;
      patterns[10466] = 33'b1010111101100010_0_0_00_000_000_000_0_0_00;
      patterns[10467] = 33'b1011011101100010_0_1_11_110_010_111_0_x_00;
      patterns[10468] = 33'b1011111101100010_1_1_11_110_010_111_0_x_00;
      patterns[10469] = 33'b1011111101100010_0_0_00_000_000_000_0_0_00;
      patterns[10470] = 33'b0101011101100000_0_1_xx_110_xxx_111_0_1_01;
      patterns[10471] = 33'b0101111101100000_1_1_xx_110_xxx_111_0_1_01;
      patterns[10472] = 33'b0101111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10473] = 33'b0100011101100000_0_0_xx_110_111_xxx_1_x_xx;
      patterns[10474] = 33'b0100111101100000_1_0_xx_110_111_xxx_1_x_xx;
      patterns[10475] = 33'b0100111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10476] = 33'b0000011101111110_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10477] = 33'b0000111101111110_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10478] = 33'b0000111101111110_0_0_00_000_000_000_0_0_00;
      patterns[10479] = 33'b1000011101100011_0_1_00_110_011_111_0_x_00;
      patterns[10480] = 33'b1000111101100011_1_1_00_110_011_111_0_x_00;
      patterns[10481] = 33'b1000111101100011_0_0_00_000_000_000_0_0_00;
      patterns[10482] = 33'b1001011101100011_0_1_01_110_011_111_0_x_00;
      patterns[10483] = 33'b1001111101100011_1_1_01_110_011_111_0_x_00;
      patterns[10484] = 33'b1001111101100011_0_0_00_000_000_000_0_0_00;
      patterns[10485] = 33'b1010011101100011_0_1_10_110_011_111_0_x_00;
      patterns[10486] = 33'b1010111101100011_1_1_10_110_011_111_0_x_00;
      patterns[10487] = 33'b1010111101100011_0_0_00_000_000_000_0_0_00;
      patterns[10488] = 33'b1011011101100011_0_1_11_110_011_111_0_x_00;
      patterns[10489] = 33'b1011111101100011_1_1_11_110_011_111_0_x_00;
      patterns[10490] = 33'b1011111101100011_0_0_00_000_000_000_0_0_00;
      patterns[10491] = 33'b0101011101100000_0_1_xx_110_xxx_111_0_1_01;
      patterns[10492] = 33'b0101111101100000_1_1_xx_110_xxx_111_0_1_01;
      patterns[10493] = 33'b0101111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10494] = 33'b0100011101100000_0_0_xx_110_111_xxx_1_x_xx;
      patterns[10495] = 33'b0100111101100000_1_0_xx_110_111_xxx_1_x_xx;
      patterns[10496] = 33'b0100111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10497] = 33'b0000011101110111_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10498] = 33'b0000111101110111_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10499] = 33'b0000111101110111_0_0_00_000_000_000_0_0_00;
      patterns[10500] = 33'b1000011101100100_0_1_00_110_100_111_0_x_00;
      patterns[10501] = 33'b1000111101100100_1_1_00_110_100_111_0_x_00;
      patterns[10502] = 33'b1000111101100100_0_0_00_000_000_000_0_0_00;
      patterns[10503] = 33'b1001011101100100_0_1_01_110_100_111_0_x_00;
      patterns[10504] = 33'b1001111101100100_1_1_01_110_100_111_0_x_00;
      patterns[10505] = 33'b1001111101100100_0_0_00_000_000_000_0_0_00;
      patterns[10506] = 33'b1010011101100100_0_1_10_110_100_111_0_x_00;
      patterns[10507] = 33'b1010111101100100_1_1_10_110_100_111_0_x_00;
      patterns[10508] = 33'b1010111101100100_0_0_00_000_000_000_0_0_00;
      patterns[10509] = 33'b1011011101100100_0_1_11_110_100_111_0_x_00;
      patterns[10510] = 33'b1011111101100100_1_1_11_110_100_111_0_x_00;
      patterns[10511] = 33'b1011111101100100_0_0_00_000_000_000_0_0_00;
      patterns[10512] = 33'b0101011101100000_0_1_xx_110_xxx_111_0_1_01;
      patterns[10513] = 33'b0101111101100000_1_1_xx_110_xxx_111_0_1_01;
      patterns[10514] = 33'b0101111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10515] = 33'b0100011101100000_0_0_xx_110_111_xxx_1_x_xx;
      patterns[10516] = 33'b0100111101100000_1_0_xx_110_111_xxx_1_x_xx;
      patterns[10517] = 33'b0100111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10518] = 33'b0000011101001100_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10519] = 33'b0000111101001100_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10520] = 33'b0000111101001100_0_0_00_000_000_000_0_0_00;
      patterns[10521] = 33'b1000011101100101_0_1_00_110_101_111_0_x_00;
      patterns[10522] = 33'b1000111101100101_1_1_00_110_101_111_0_x_00;
      patterns[10523] = 33'b1000111101100101_0_0_00_000_000_000_0_0_00;
      patterns[10524] = 33'b1001011101100101_0_1_01_110_101_111_0_x_00;
      patterns[10525] = 33'b1001111101100101_1_1_01_110_101_111_0_x_00;
      patterns[10526] = 33'b1001111101100101_0_0_00_000_000_000_0_0_00;
      patterns[10527] = 33'b1010011101100101_0_1_10_110_101_111_0_x_00;
      patterns[10528] = 33'b1010111101100101_1_1_10_110_101_111_0_x_00;
      patterns[10529] = 33'b1010111101100101_0_0_00_000_000_000_0_0_00;
      patterns[10530] = 33'b1011011101100101_0_1_11_110_101_111_0_x_00;
      patterns[10531] = 33'b1011111101100101_1_1_11_110_101_111_0_x_00;
      patterns[10532] = 33'b1011111101100101_0_0_00_000_000_000_0_0_00;
      patterns[10533] = 33'b0101011101100000_0_1_xx_110_xxx_111_0_1_01;
      patterns[10534] = 33'b0101111101100000_1_1_xx_110_xxx_111_0_1_01;
      patterns[10535] = 33'b0101111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10536] = 33'b0100011101100000_0_0_xx_110_111_xxx_1_x_xx;
      patterns[10537] = 33'b0100111101100000_1_0_xx_110_111_xxx_1_x_xx;
      patterns[10538] = 33'b0100111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10539] = 33'b0000011101011011_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10540] = 33'b0000111101011011_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10541] = 33'b0000111101011011_0_0_00_000_000_000_0_0_00;
      patterns[10542] = 33'b1000011101100110_0_1_00_110_110_111_0_x_00;
      patterns[10543] = 33'b1000111101100110_1_1_00_110_110_111_0_x_00;
      patterns[10544] = 33'b1000111101100110_0_0_00_000_000_000_0_0_00;
      patterns[10545] = 33'b1001011101100110_0_1_01_110_110_111_0_x_00;
      patterns[10546] = 33'b1001111101100110_1_1_01_110_110_111_0_x_00;
      patterns[10547] = 33'b1001111101100110_0_0_00_000_000_000_0_0_00;
      patterns[10548] = 33'b1010011101100110_0_1_10_110_110_111_0_x_00;
      patterns[10549] = 33'b1010111101100110_1_1_10_110_110_111_0_x_00;
      patterns[10550] = 33'b1010111101100110_0_0_00_000_000_000_0_0_00;
      patterns[10551] = 33'b1011011101100110_0_1_11_110_110_111_0_x_00;
      patterns[10552] = 33'b1011111101100110_1_1_11_110_110_111_0_x_00;
      patterns[10553] = 33'b1011111101100110_0_0_00_000_000_000_0_0_00;
      patterns[10554] = 33'b0101011101100000_0_1_xx_110_xxx_111_0_1_01;
      patterns[10555] = 33'b0101111101100000_1_1_xx_110_xxx_111_0_1_01;
      patterns[10556] = 33'b0101111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10557] = 33'b0100011101100000_0_0_xx_110_111_xxx_1_x_xx;
      patterns[10558] = 33'b0100111101100000_1_0_xx_110_111_xxx_1_x_xx;
      patterns[10559] = 33'b0100111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10560] = 33'b0000011110100101_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10561] = 33'b0000111110100101_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10562] = 33'b0000111110100101_0_0_00_000_000_000_0_0_00;
      patterns[10563] = 33'b1000011101100111_0_1_00_110_111_111_0_x_00;
      patterns[10564] = 33'b1000111101100111_1_1_00_110_111_111_0_x_00;
      patterns[10565] = 33'b1000111101100111_0_0_00_000_000_000_0_0_00;
      patterns[10566] = 33'b1001011101100111_0_1_01_110_111_111_0_x_00;
      patterns[10567] = 33'b1001111101100111_1_1_01_110_111_111_0_x_00;
      patterns[10568] = 33'b1001111101100111_0_0_00_000_000_000_0_0_00;
      patterns[10569] = 33'b1010011101100111_0_1_10_110_111_111_0_x_00;
      patterns[10570] = 33'b1010111101100111_1_1_10_110_111_111_0_x_00;
      patterns[10571] = 33'b1010111101100111_0_0_00_000_000_000_0_0_00;
      patterns[10572] = 33'b1011011101100111_0_1_11_110_111_111_0_x_00;
      patterns[10573] = 33'b1011111101100111_1_1_11_110_111_111_0_x_00;
      patterns[10574] = 33'b1011111101100111_0_0_00_000_000_000_0_0_00;
      patterns[10575] = 33'b0101011101100000_0_1_xx_110_xxx_111_0_1_01;
      patterns[10576] = 33'b0101111101100000_1_1_xx_110_xxx_111_0_1_01;
      patterns[10577] = 33'b0101111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10578] = 33'b0100011101100000_0_0_xx_110_111_xxx_1_x_xx;
      patterns[10579] = 33'b0100111101100000_1_0_xx_110_111_xxx_1_x_xx;
      patterns[10580] = 33'b0100111101100000_0_0_00_000_000_000_0_0_00;
      patterns[10581] = 33'b0000011110001100_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10582] = 33'b0000111110001100_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10583] = 33'b0000111110001100_0_0_00_000_000_000_0_0_00;
      patterns[10584] = 33'b1000011101110000_0_1_00_111_000_111_0_x_00;
      patterns[10585] = 33'b1000111101110000_1_1_00_111_000_111_0_x_00;
      patterns[10586] = 33'b1000111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10587] = 33'b1001011101110000_0_1_01_111_000_111_0_x_00;
      patterns[10588] = 33'b1001111101110000_1_1_01_111_000_111_0_x_00;
      patterns[10589] = 33'b1001111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10590] = 33'b1010011101110000_0_1_10_111_000_111_0_x_00;
      patterns[10591] = 33'b1010111101110000_1_1_10_111_000_111_0_x_00;
      patterns[10592] = 33'b1010111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10593] = 33'b1011011101110000_0_1_11_111_000_111_0_x_00;
      patterns[10594] = 33'b1011111101110000_1_1_11_111_000_111_0_x_00;
      patterns[10595] = 33'b1011111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10596] = 33'b0101011101110000_0_1_xx_111_xxx_111_0_1_01;
      patterns[10597] = 33'b0101111101110000_1_1_xx_111_xxx_111_0_1_01;
      patterns[10598] = 33'b0101111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10599] = 33'b0100011101110000_0_0_xx_111_111_xxx_1_x_xx;
      patterns[10600] = 33'b0100111101110000_1_0_xx_111_111_xxx_1_x_xx;
      patterns[10601] = 33'b0100111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10602] = 33'b0000011100111011_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10603] = 33'b0000111100111011_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10604] = 33'b0000111100111011_0_0_00_000_000_000_0_0_00;
      patterns[10605] = 33'b1000011101110001_0_1_00_111_001_111_0_x_00;
      patterns[10606] = 33'b1000111101110001_1_1_00_111_001_111_0_x_00;
      patterns[10607] = 33'b1000111101110001_0_0_00_000_000_000_0_0_00;
      patterns[10608] = 33'b1001011101110001_0_1_01_111_001_111_0_x_00;
      patterns[10609] = 33'b1001111101110001_1_1_01_111_001_111_0_x_00;
      patterns[10610] = 33'b1001111101110001_0_0_00_000_000_000_0_0_00;
      patterns[10611] = 33'b1010011101110001_0_1_10_111_001_111_0_x_00;
      patterns[10612] = 33'b1010111101110001_1_1_10_111_001_111_0_x_00;
      patterns[10613] = 33'b1010111101110001_0_0_00_000_000_000_0_0_00;
      patterns[10614] = 33'b1011011101110001_0_1_11_111_001_111_0_x_00;
      patterns[10615] = 33'b1011111101110001_1_1_11_111_001_111_0_x_00;
      patterns[10616] = 33'b1011111101110001_0_0_00_000_000_000_0_0_00;
      patterns[10617] = 33'b0101011101110000_0_1_xx_111_xxx_111_0_1_01;
      patterns[10618] = 33'b0101111101110000_1_1_xx_111_xxx_111_0_1_01;
      patterns[10619] = 33'b0101111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10620] = 33'b0100011101110000_0_0_xx_111_111_xxx_1_x_xx;
      patterns[10621] = 33'b0100111101110000_1_0_xx_111_111_xxx_1_x_xx;
      patterns[10622] = 33'b0100111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10623] = 33'b0000011101001000_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10624] = 33'b0000111101001000_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10625] = 33'b0000111101001000_0_0_00_000_000_000_0_0_00;
      patterns[10626] = 33'b1000011101110010_0_1_00_111_010_111_0_x_00;
      patterns[10627] = 33'b1000111101110010_1_1_00_111_010_111_0_x_00;
      patterns[10628] = 33'b1000111101110010_0_0_00_000_000_000_0_0_00;
      patterns[10629] = 33'b1001011101110010_0_1_01_111_010_111_0_x_00;
      patterns[10630] = 33'b1001111101110010_1_1_01_111_010_111_0_x_00;
      patterns[10631] = 33'b1001111101110010_0_0_00_000_000_000_0_0_00;
      patterns[10632] = 33'b1010011101110010_0_1_10_111_010_111_0_x_00;
      patterns[10633] = 33'b1010111101110010_1_1_10_111_010_111_0_x_00;
      patterns[10634] = 33'b1010111101110010_0_0_00_000_000_000_0_0_00;
      patterns[10635] = 33'b1011011101110010_0_1_11_111_010_111_0_x_00;
      patterns[10636] = 33'b1011111101110010_1_1_11_111_010_111_0_x_00;
      patterns[10637] = 33'b1011111101110010_0_0_00_000_000_000_0_0_00;
      patterns[10638] = 33'b0101011101110000_0_1_xx_111_xxx_111_0_1_01;
      patterns[10639] = 33'b0101111101110000_1_1_xx_111_xxx_111_0_1_01;
      patterns[10640] = 33'b0101111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10641] = 33'b0100011101110000_0_0_xx_111_111_xxx_1_x_xx;
      patterns[10642] = 33'b0100111101110000_1_0_xx_111_111_xxx_1_x_xx;
      patterns[10643] = 33'b0100111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10644] = 33'b0000011111011000_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10645] = 33'b0000111111011000_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10646] = 33'b0000111111011000_0_0_00_000_000_000_0_0_00;
      patterns[10647] = 33'b1000011101110011_0_1_00_111_011_111_0_x_00;
      patterns[10648] = 33'b1000111101110011_1_1_00_111_011_111_0_x_00;
      patterns[10649] = 33'b1000111101110011_0_0_00_000_000_000_0_0_00;
      patterns[10650] = 33'b1001011101110011_0_1_01_111_011_111_0_x_00;
      patterns[10651] = 33'b1001111101110011_1_1_01_111_011_111_0_x_00;
      patterns[10652] = 33'b1001111101110011_0_0_00_000_000_000_0_0_00;
      patterns[10653] = 33'b1010011101110011_0_1_10_111_011_111_0_x_00;
      patterns[10654] = 33'b1010111101110011_1_1_10_111_011_111_0_x_00;
      patterns[10655] = 33'b1010111101110011_0_0_00_000_000_000_0_0_00;
      patterns[10656] = 33'b1011011101110011_0_1_11_111_011_111_0_x_00;
      patterns[10657] = 33'b1011111101110011_1_1_11_111_011_111_0_x_00;
      patterns[10658] = 33'b1011111101110011_0_0_00_000_000_000_0_0_00;
      patterns[10659] = 33'b0101011101110000_0_1_xx_111_xxx_111_0_1_01;
      patterns[10660] = 33'b0101111101110000_1_1_xx_111_xxx_111_0_1_01;
      patterns[10661] = 33'b0101111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10662] = 33'b0100011101110000_0_0_xx_111_111_xxx_1_x_xx;
      patterns[10663] = 33'b0100111101110000_1_0_xx_111_111_xxx_1_x_xx;
      patterns[10664] = 33'b0100111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10665] = 33'b0000011100011101_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10666] = 33'b0000111100011101_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10667] = 33'b0000111100011101_0_0_00_000_000_000_0_0_00;
      patterns[10668] = 33'b1000011101110100_0_1_00_111_100_111_0_x_00;
      patterns[10669] = 33'b1000111101110100_1_1_00_111_100_111_0_x_00;
      patterns[10670] = 33'b1000111101110100_0_0_00_000_000_000_0_0_00;
      patterns[10671] = 33'b1001011101110100_0_1_01_111_100_111_0_x_00;
      patterns[10672] = 33'b1001111101110100_1_1_01_111_100_111_0_x_00;
      patterns[10673] = 33'b1001111101110100_0_0_00_000_000_000_0_0_00;
      patterns[10674] = 33'b1010011101110100_0_1_10_111_100_111_0_x_00;
      patterns[10675] = 33'b1010111101110100_1_1_10_111_100_111_0_x_00;
      patterns[10676] = 33'b1010111101110100_0_0_00_000_000_000_0_0_00;
      patterns[10677] = 33'b1011011101110100_0_1_11_111_100_111_0_x_00;
      patterns[10678] = 33'b1011111101110100_1_1_11_111_100_111_0_x_00;
      patterns[10679] = 33'b1011111101110100_0_0_00_000_000_000_0_0_00;
      patterns[10680] = 33'b0101011101110000_0_1_xx_111_xxx_111_0_1_01;
      patterns[10681] = 33'b0101111101110000_1_1_xx_111_xxx_111_0_1_01;
      patterns[10682] = 33'b0101111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10683] = 33'b0100011101110000_0_0_xx_111_111_xxx_1_x_xx;
      patterns[10684] = 33'b0100111101110000_1_0_xx_111_111_xxx_1_x_xx;
      patterns[10685] = 33'b0100111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10686] = 33'b0000011101011010_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10687] = 33'b0000111101011010_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10688] = 33'b0000111101011010_0_0_00_000_000_000_0_0_00;
      patterns[10689] = 33'b1000011101110101_0_1_00_111_101_111_0_x_00;
      patterns[10690] = 33'b1000111101110101_1_1_00_111_101_111_0_x_00;
      patterns[10691] = 33'b1000111101110101_0_0_00_000_000_000_0_0_00;
      patterns[10692] = 33'b1001011101110101_0_1_01_111_101_111_0_x_00;
      patterns[10693] = 33'b1001111101110101_1_1_01_111_101_111_0_x_00;
      patterns[10694] = 33'b1001111101110101_0_0_00_000_000_000_0_0_00;
      patterns[10695] = 33'b1010011101110101_0_1_10_111_101_111_0_x_00;
      patterns[10696] = 33'b1010111101110101_1_1_10_111_101_111_0_x_00;
      patterns[10697] = 33'b1010111101110101_0_0_00_000_000_000_0_0_00;
      patterns[10698] = 33'b1011011101110101_0_1_11_111_101_111_0_x_00;
      patterns[10699] = 33'b1011111101110101_1_1_11_111_101_111_0_x_00;
      patterns[10700] = 33'b1011111101110101_0_0_00_000_000_000_0_0_00;
      patterns[10701] = 33'b0101011101110000_0_1_xx_111_xxx_111_0_1_01;
      patterns[10702] = 33'b0101111101110000_1_1_xx_111_xxx_111_0_1_01;
      patterns[10703] = 33'b0101111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10704] = 33'b0100011101110000_0_0_xx_111_111_xxx_1_x_xx;
      patterns[10705] = 33'b0100111101110000_1_0_xx_111_111_xxx_1_x_xx;
      patterns[10706] = 33'b0100111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10707] = 33'b0000011100001110_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10708] = 33'b0000111100001110_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10709] = 33'b0000111100001110_0_0_00_000_000_000_0_0_00;
      patterns[10710] = 33'b1000011101110110_0_1_00_111_110_111_0_x_00;
      patterns[10711] = 33'b1000111101110110_1_1_00_111_110_111_0_x_00;
      patterns[10712] = 33'b1000111101110110_0_0_00_000_000_000_0_0_00;
      patterns[10713] = 33'b1001011101110110_0_1_01_111_110_111_0_x_00;
      patterns[10714] = 33'b1001111101110110_1_1_01_111_110_111_0_x_00;
      patterns[10715] = 33'b1001111101110110_0_0_00_000_000_000_0_0_00;
      patterns[10716] = 33'b1010011101110110_0_1_10_111_110_111_0_x_00;
      patterns[10717] = 33'b1010111101110110_1_1_10_111_110_111_0_x_00;
      patterns[10718] = 33'b1010111101110110_0_0_00_000_000_000_0_0_00;
      patterns[10719] = 33'b1011011101110110_0_1_11_111_110_111_0_x_00;
      patterns[10720] = 33'b1011111101110110_1_1_11_111_110_111_0_x_00;
      patterns[10721] = 33'b1011111101110110_0_0_00_000_000_000_0_0_00;
      patterns[10722] = 33'b0101011101110000_0_1_xx_111_xxx_111_0_1_01;
      patterns[10723] = 33'b0101111101110000_1_1_xx_111_xxx_111_0_1_01;
      patterns[10724] = 33'b0101111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10725] = 33'b0100011101110000_0_0_xx_111_111_xxx_1_x_xx;
      patterns[10726] = 33'b0100111101110000_1_0_xx_111_111_xxx_1_x_xx;
      patterns[10727] = 33'b0100111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10728] = 33'b0000011101000011_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10729] = 33'b0000111101000011_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10730] = 33'b0000111101000011_0_0_00_000_000_000_0_0_00;
      patterns[10731] = 33'b1000011101110111_0_1_00_111_111_111_0_x_00;
      patterns[10732] = 33'b1000111101110111_1_1_00_111_111_111_0_x_00;
      patterns[10733] = 33'b1000111101110111_0_0_00_000_000_000_0_0_00;
      patterns[10734] = 33'b1001011101110111_0_1_01_111_111_111_0_x_00;
      patterns[10735] = 33'b1001111101110111_1_1_01_111_111_111_0_x_00;
      patterns[10736] = 33'b1001111101110111_0_0_00_000_000_000_0_0_00;
      patterns[10737] = 33'b1010011101110111_0_1_10_111_111_111_0_x_00;
      patterns[10738] = 33'b1010111101110111_1_1_10_111_111_111_0_x_00;
      patterns[10739] = 33'b1010111101110111_0_0_00_000_000_000_0_0_00;
      patterns[10740] = 33'b1011011101110111_0_1_11_111_111_111_0_x_00;
      patterns[10741] = 33'b1011111101110111_1_1_11_111_111_111_0_x_00;
      patterns[10742] = 33'b1011111101110111_0_0_00_000_000_000_0_0_00;
      patterns[10743] = 33'b0101011101110000_0_1_xx_111_xxx_111_0_1_01;
      patterns[10744] = 33'b0101111101110000_1_1_xx_111_xxx_111_0_1_01;
      patterns[10745] = 33'b0101111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10746] = 33'b0100011101110000_0_0_xx_111_111_xxx_1_x_xx;
      patterns[10747] = 33'b0100111101110000_1_0_xx_111_111_xxx_1_x_xx;
      patterns[10748] = 33'b0100111101110000_0_0_00_000_000_000_0_0_00;
      patterns[10749] = 33'b0000011101100010_0_1_xx_xxx_xxx_111_0_x_10;
      patterns[10750] = 33'b0000111101100010_1_1_xx_xxx_xxx_111_0_x_10;
      patterns[10751] = 33'b0000111101100010_0_0_00_000_000_000_0_0_00;

      for (i = 0; i < 10752; i = i + 1)
      begin
        INST = patterns[i][32:17];
        FL_Z = patterns[i][16];
        #10;
        if (patterns[i][15] !== 1'hx)
        begin
          if (WE !== patterns[i][15])
          begin
            $display("%d:WE: (assertion error). Expected %h, found %h", i, patterns[i][15], WE);
            $finish;
          end
        end
        if (patterns[i][14:13] !== 2'hx)
        begin
          if (ALUOP !== patterns[i][14:13])
          begin
            $display("%d:ALUOP: (assertion error). Expected %h, found %h", i, patterns[i][14:13], ALUOP);
            $finish;
          end
        end
        if (patterns[i][12:10] !== 3'hx)
        begin
          if (RS1 !== patterns[i][12:10])
          begin
            $display("%d:RS1: (assertion error). Expected %h, found %h", i, patterns[i][12:10], RS1);
            $finish;
          end
        end
        if (patterns[i][9:7] !== 3'hx)
        begin
          if (RS2 !== patterns[i][9:7])
          begin
            $display("%d:RS2: (assertion error). Expected %h, found %h", i, patterns[i][9:7], RS2);
            $finish;
          end
        end
        if (patterns[i][6:4] !== 3'hx)
        begin
          if (WS !== patterns[i][6:4])
          begin
            $display("%d:WS: (assertion error). Expected %h, found %h", i, patterns[i][6:4], WS);
            $finish;
          end
        end
        if (patterns[i][3] !== 1'hx)
        begin
          if (STR !== patterns[i][3])
          begin
            $display("%d:STR: (assertion error). Expected %h, found %h", i, patterns[i][3], STR);
            $finish;
          end
        end
        if (patterns[i][2] !== 1'hx)
        begin
          if (LDR !== patterns[i][2])
          begin
            $display("%d:LDR: (assertion error). Expected %h, found %h", i, patterns[i][2], LDR);
            $finish;
          end
        end
        if (patterns[i][1:0] !== 2'hx)
        begin
          if (DMUX !== patterns[i][1:0])
          begin
            $display("%d:DMUX: (assertion error). Expected %h, found %h", i, patterns[i][1:0], DMUX);
            $finish;
          end
        end
      end

      $display("All tests passed.");
    end
    endmodule
