--  A testbench for control_unit_RS1_tb
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity control_unit_RS1_tb is
end control_unit_RS1_tb;

architecture behav of control_unit_RS1_tb is
  component main
    port (
      INST: in std_logic_vector(15 downto 0);
      ALUOP: out std_logic_vector(1 downto 0);
      RS1: out std_logic_vector(2 downto 0);
      RS2: out std_logic_vector(2 downto 0);
      WS: out std_logic_vector(2 downto 0);
      STR: out std_logic;
      WE: out std_logic;
      DMUX: out std_logic_vector(1 downto 0);
      LDR: out std_logic);
  end component;

  signal INST : std_logic_vector(15 downto 0);
  signal ALUOP : std_logic_vector(1 downto 0);
  signal RS1 : std_logic_vector(2 downto 0);
  signal RS2 : std_logic_vector(2 downto 0);
  signal WS : std_logic_vector(2 downto 0);
  signal STR : std_logic;
  signal WE : std_logic;
  signal DMUX : std_logic_vector(1 downto 0);
  signal LDR : std_logic;
  function to_string ( a: std_logic_vector) return string is
      variable b : string (1 to a'length) := (others => NUL);
      variable stri : integer := 1; 
  begin
      for i in a'range loop
          b(stri) := std_logic'image(a((i)))(2);
      stri := stri+1;
      end loop;
      return b;
  end function;
begin
  main_0 : main port map (
    INST => INST,
    ALUOP => ALUOP,
    RS1 => RS1,
    RS2 => RS2,
    WS => WS,
    STR => STR,
    WE => WE,
    DMUX => DMUX,
    LDR => LDR );
  process
    type pattern_type is record
      INST : std_logic_vector(15 downto 0);
      RS1 : std_logic_vector(2 downto 0);
    end record;
    type pattern_array is array (natural range <>) of pattern_type;
    constant patterns : pattern_array := (
      ("1000000000000000", "000"), -- i=0
      ("1001000000000000", "000"), -- i=1
      ("1010000000000000", "000"), -- i=2
      ("1011000000000000", "000"), -- i=3
      ("0101000000000000", "000"), -- i=4
      ("0100000000000000", "000"), -- i=5
      ("1000000000000001", "000"), -- i=6
      ("1001000000000001", "000"), -- i=7
      ("1010000000000001", "000"), -- i=8
      ("1011000000000001", "000"), -- i=9
      ("0101000000000000", "000"), -- i=10
      ("0100000000000000", "000"), -- i=11
      ("1000000000000010", "000"), -- i=12
      ("1001000000000010", "000"), -- i=13
      ("1010000000000010", "000"), -- i=14
      ("1011000000000010", "000"), -- i=15
      ("0101000000000000", "000"), -- i=16
      ("0100000000000000", "000"), -- i=17
      ("1000000000000011", "000"), -- i=18
      ("1001000000000011", "000"), -- i=19
      ("1010000000000011", "000"), -- i=20
      ("1011000000000011", "000"), -- i=21
      ("0101000000000000", "000"), -- i=22
      ("0100000000000000", "000"), -- i=23
      ("1000000000000100", "000"), -- i=24
      ("1001000000000100", "000"), -- i=25
      ("1010000000000100", "000"), -- i=26
      ("1011000000000100", "000"), -- i=27
      ("0101000000000000", "000"), -- i=28
      ("0100000000000000", "000"), -- i=29
      ("1000000000000101", "000"), -- i=30
      ("1001000000000101", "000"), -- i=31
      ("1010000000000101", "000"), -- i=32
      ("1011000000000101", "000"), -- i=33
      ("0101000000000000", "000"), -- i=34
      ("0100000000000000", "000"), -- i=35
      ("1000000000000110", "000"), -- i=36
      ("1001000000000110", "000"), -- i=37
      ("1010000000000110", "000"), -- i=38
      ("1011000000000110", "000"), -- i=39
      ("0101000000000000", "000"), -- i=40
      ("0100000000000000", "000"), -- i=41
      ("1000000000000111", "000"), -- i=42
      ("1001000000000111", "000"), -- i=43
      ("1010000000000111", "000"), -- i=44
      ("1011000000000111", "000"), -- i=45
      ("0101000000000000", "000"), -- i=46
      ("0100000000000000", "000"), -- i=47
      ("1000000000010000", "001"), -- i=48
      ("1001000000010000", "001"), -- i=49
      ("1010000000010000", "001"), -- i=50
      ("1011000000010000", "001"), -- i=51
      ("0101000000010000", "001"), -- i=52
      ("0100000000010000", "001"), -- i=53
      ("1000000000010001", "001"), -- i=54
      ("1001000000010001", "001"), -- i=55
      ("1010000000010001", "001"), -- i=56
      ("1011000000010001", "001"), -- i=57
      ("0101000000010000", "001"), -- i=58
      ("0100000000010000", "001"), -- i=59
      ("1000000000010010", "001"), -- i=60
      ("1001000000010010", "001"), -- i=61
      ("1010000000010010", "001"), -- i=62
      ("1011000000010010", "001"), -- i=63
      ("0101000000010000", "001"), -- i=64
      ("0100000000010000", "001"), -- i=65
      ("1000000000010011", "001"), -- i=66
      ("1001000000010011", "001"), -- i=67
      ("1010000000010011", "001"), -- i=68
      ("1011000000010011", "001"), -- i=69
      ("0101000000010000", "001"), -- i=70
      ("0100000000010000", "001"), -- i=71
      ("1000000000010100", "001"), -- i=72
      ("1001000000010100", "001"), -- i=73
      ("1010000000010100", "001"), -- i=74
      ("1011000000010100", "001"), -- i=75
      ("0101000000010000", "001"), -- i=76
      ("0100000000010000", "001"), -- i=77
      ("1000000000010101", "001"), -- i=78
      ("1001000000010101", "001"), -- i=79
      ("1010000000010101", "001"), -- i=80
      ("1011000000010101", "001"), -- i=81
      ("0101000000010000", "001"), -- i=82
      ("0100000000010000", "001"), -- i=83
      ("1000000000010110", "001"), -- i=84
      ("1001000000010110", "001"), -- i=85
      ("1010000000010110", "001"), -- i=86
      ("1011000000010110", "001"), -- i=87
      ("0101000000010000", "001"), -- i=88
      ("0100000000010000", "001"), -- i=89
      ("1000000000010111", "001"), -- i=90
      ("1001000000010111", "001"), -- i=91
      ("1010000000010111", "001"), -- i=92
      ("1011000000010111", "001"), -- i=93
      ("0101000000010000", "001"), -- i=94
      ("0100000000010000", "001"), -- i=95
      ("1000000000100000", "010"), -- i=96
      ("1001000000100000", "010"), -- i=97
      ("1010000000100000", "010"), -- i=98
      ("1011000000100000", "010"), -- i=99
      ("0101000000100000", "010"), -- i=100
      ("0100000000100000", "010"), -- i=101
      ("1000000000100001", "010"), -- i=102
      ("1001000000100001", "010"), -- i=103
      ("1010000000100001", "010"), -- i=104
      ("1011000000100001", "010"), -- i=105
      ("0101000000100000", "010"), -- i=106
      ("0100000000100000", "010"), -- i=107
      ("1000000000100010", "010"), -- i=108
      ("1001000000100010", "010"), -- i=109
      ("1010000000100010", "010"), -- i=110
      ("1011000000100010", "010"), -- i=111
      ("0101000000100000", "010"), -- i=112
      ("0100000000100000", "010"), -- i=113
      ("1000000000100011", "010"), -- i=114
      ("1001000000100011", "010"), -- i=115
      ("1010000000100011", "010"), -- i=116
      ("1011000000100011", "010"), -- i=117
      ("0101000000100000", "010"), -- i=118
      ("0100000000100000", "010"), -- i=119
      ("1000000000100100", "010"), -- i=120
      ("1001000000100100", "010"), -- i=121
      ("1010000000100100", "010"), -- i=122
      ("1011000000100100", "010"), -- i=123
      ("0101000000100000", "010"), -- i=124
      ("0100000000100000", "010"), -- i=125
      ("1000000000100101", "010"), -- i=126
      ("1001000000100101", "010"), -- i=127
      ("1010000000100101", "010"), -- i=128
      ("1011000000100101", "010"), -- i=129
      ("0101000000100000", "010"), -- i=130
      ("0100000000100000", "010"), -- i=131
      ("1000000000100110", "010"), -- i=132
      ("1001000000100110", "010"), -- i=133
      ("1010000000100110", "010"), -- i=134
      ("1011000000100110", "010"), -- i=135
      ("0101000000100000", "010"), -- i=136
      ("0100000000100000", "010"), -- i=137
      ("1000000000100111", "010"), -- i=138
      ("1001000000100111", "010"), -- i=139
      ("1010000000100111", "010"), -- i=140
      ("1011000000100111", "010"), -- i=141
      ("0101000000100000", "010"), -- i=142
      ("0100000000100000", "010"), -- i=143
      ("1000000000110000", "011"), -- i=144
      ("1001000000110000", "011"), -- i=145
      ("1010000000110000", "011"), -- i=146
      ("1011000000110000", "011"), -- i=147
      ("0101000000110000", "011"), -- i=148
      ("0100000000110000", "011"), -- i=149
      ("1000000000110001", "011"), -- i=150
      ("1001000000110001", "011"), -- i=151
      ("1010000000110001", "011"), -- i=152
      ("1011000000110001", "011"), -- i=153
      ("0101000000110000", "011"), -- i=154
      ("0100000000110000", "011"), -- i=155
      ("1000000000110010", "011"), -- i=156
      ("1001000000110010", "011"), -- i=157
      ("1010000000110010", "011"), -- i=158
      ("1011000000110010", "011"), -- i=159
      ("0101000000110000", "011"), -- i=160
      ("0100000000110000", "011"), -- i=161
      ("1000000000110011", "011"), -- i=162
      ("1001000000110011", "011"), -- i=163
      ("1010000000110011", "011"), -- i=164
      ("1011000000110011", "011"), -- i=165
      ("0101000000110000", "011"), -- i=166
      ("0100000000110000", "011"), -- i=167
      ("1000000000110100", "011"), -- i=168
      ("1001000000110100", "011"), -- i=169
      ("1010000000110100", "011"), -- i=170
      ("1011000000110100", "011"), -- i=171
      ("0101000000110000", "011"), -- i=172
      ("0100000000110000", "011"), -- i=173
      ("1000000000110101", "011"), -- i=174
      ("1001000000110101", "011"), -- i=175
      ("1010000000110101", "011"), -- i=176
      ("1011000000110101", "011"), -- i=177
      ("0101000000110000", "011"), -- i=178
      ("0100000000110000", "011"), -- i=179
      ("1000000000110110", "011"), -- i=180
      ("1001000000110110", "011"), -- i=181
      ("1010000000110110", "011"), -- i=182
      ("1011000000110110", "011"), -- i=183
      ("0101000000110000", "011"), -- i=184
      ("0100000000110000", "011"), -- i=185
      ("1000000000110111", "011"), -- i=186
      ("1001000000110111", "011"), -- i=187
      ("1010000000110111", "011"), -- i=188
      ("1011000000110111", "011"), -- i=189
      ("0101000000110000", "011"), -- i=190
      ("0100000000110000", "011"), -- i=191
      ("1000000001000000", "100"), -- i=192
      ("1001000001000000", "100"), -- i=193
      ("1010000001000000", "100"), -- i=194
      ("1011000001000000", "100"), -- i=195
      ("0101000001000000", "100"), -- i=196
      ("0100000001000000", "100"), -- i=197
      ("1000000001000001", "100"), -- i=198
      ("1001000001000001", "100"), -- i=199
      ("1010000001000001", "100"), -- i=200
      ("1011000001000001", "100"), -- i=201
      ("0101000001000000", "100"), -- i=202
      ("0100000001000000", "100"), -- i=203
      ("1000000001000010", "100"), -- i=204
      ("1001000001000010", "100"), -- i=205
      ("1010000001000010", "100"), -- i=206
      ("1011000001000010", "100"), -- i=207
      ("0101000001000000", "100"), -- i=208
      ("0100000001000000", "100"), -- i=209
      ("1000000001000011", "100"), -- i=210
      ("1001000001000011", "100"), -- i=211
      ("1010000001000011", "100"), -- i=212
      ("1011000001000011", "100"), -- i=213
      ("0101000001000000", "100"), -- i=214
      ("0100000001000000", "100"), -- i=215
      ("1000000001000100", "100"), -- i=216
      ("1001000001000100", "100"), -- i=217
      ("1010000001000100", "100"), -- i=218
      ("1011000001000100", "100"), -- i=219
      ("0101000001000000", "100"), -- i=220
      ("0100000001000000", "100"), -- i=221
      ("1000000001000101", "100"), -- i=222
      ("1001000001000101", "100"), -- i=223
      ("1010000001000101", "100"), -- i=224
      ("1011000001000101", "100"), -- i=225
      ("0101000001000000", "100"), -- i=226
      ("0100000001000000", "100"), -- i=227
      ("1000000001000110", "100"), -- i=228
      ("1001000001000110", "100"), -- i=229
      ("1010000001000110", "100"), -- i=230
      ("1011000001000110", "100"), -- i=231
      ("0101000001000000", "100"), -- i=232
      ("0100000001000000", "100"), -- i=233
      ("1000000001000111", "100"), -- i=234
      ("1001000001000111", "100"), -- i=235
      ("1010000001000111", "100"), -- i=236
      ("1011000001000111", "100"), -- i=237
      ("0101000001000000", "100"), -- i=238
      ("0100000001000000", "100"), -- i=239
      ("1000000001010000", "101"), -- i=240
      ("1001000001010000", "101"), -- i=241
      ("1010000001010000", "101"), -- i=242
      ("1011000001010000", "101"), -- i=243
      ("0101000001010000", "101"), -- i=244
      ("0100000001010000", "101"), -- i=245
      ("1000000001010001", "101"), -- i=246
      ("1001000001010001", "101"), -- i=247
      ("1010000001010001", "101"), -- i=248
      ("1011000001010001", "101"), -- i=249
      ("0101000001010000", "101"), -- i=250
      ("0100000001010000", "101"), -- i=251
      ("1000000001010010", "101"), -- i=252
      ("1001000001010010", "101"), -- i=253
      ("1010000001010010", "101"), -- i=254
      ("1011000001010010", "101"), -- i=255
      ("0101000001010000", "101"), -- i=256
      ("0100000001010000", "101"), -- i=257
      ("1000000001010011", "101"), -- i=258
      ("1001000001010011", "101"), -- i=259
      ("1010000001010011", "101"), -- i=260
      ("1011000001010011", "101"), -- i=261
      ("0101000001010000", "101"), -- i=262
      ("0100000001010000", "101"), -- i=263
      ("1000000001010100", "101"), -- i=264
      ("1001000001010100", "101"), -- i=265
      ("1010000001010100", "101"), -- i=266
      ("1011000001010100", "101"), -- i=267
      ("0101000001010000", "101"), -- i=268
      ("0100000001010000", "101"), -- i=269
      ("1000000001010101", "101"), -- i=270
      ("1001000001010101", "101"), -- i=271
      ("1010000001010101", "101"), -- i=272
      ("1011000001010101", "101"), -- i=273
      ("0101000001010000", "101"), -- i=274
      ("0100000001010000", "101"), -- i=275
      ("1000000001010110", "101"), -- i=276
      ("1001000001010110", "101"), -- i=277
      ("1010000001010110", "101"), -- i=278
      ("1011000001010110", "101"), -- i=279
      ("0101000001010000", "101"), -- i=280
      ("0100000001010000", "101"), -- i=281
      ("1000000001010111", "101"), -- i=282
      ("1001000001010111", "101"), -- i=283
      ("1010000001010111", "101"), -- i=284
      ("1011000001010111", "101"), -- i=285
      ("0101000001010000", "101"), -- i=286
      ("0100000001010000", "101"), -- i=287
      ("1000000001100000", "110"), -- i=288
      ("1001000001100000", "110"), -- i=289
      ("1010000001100000", "110"), -- i=290
      ("1011000001100000", "110"), -- i=291
      ("0101000001100000", "110"), -- i=292
      ("0100000001100000", "110"), -- i=293
      ("1000000001100001", "110"), -- i=294
      ("1001000001100001", "110"), -- i=295
      ("1010000001100001", "110"), -- i=296
      ("1011000001100001", "110"), -- i=297
      ("0101000001100000", "110"), -- i=298
      ("0100000001100000", "110"), -- i=299
      ("1000000001100010", "110"), -- i=300
      ("1001000001100010", "110"), -- i=301
      ("1010000001100010", "110"), -- i=302
      ("1011000001100010", "110"), -- i=303
      ("0101000001100000", "110"), -- i=304
      ("0100000001100000", "110"), -- i=305
      ("1000000001100011", "110"), -- i=306
      ("1001000001100011", "110"), -- i=307
      ("1010000001100011", "110"), -- i=308
      ("1011000001100011", "110"), -- i=309
      ("0101000001100000", "110"), -- i=310
      ("0100000001100000", "110"), -- i=311
      ("1000000001100100", "110"), -- i=312
      ("1001000001100100", "110"), -- i=313
      ("1010000001100100", "110"), -- i=314
      ("1011000001100100", "110"), -- i=315
      ("0101000001100000", "110"), -- i=316
      ("0100000001100000", "110"), -- i=317
      ("1000000001100101", "110"), -- i=318
      ("1001000001100101", "110"), -- i=319
      ("1010000001100101", "110"), -- i=320
      ("1011000001100101", "110"), -- i=321
      ("0101000001100000", "110"), -- i=322
      ("0100000001100000", "110"), -- i=323
      ("1000000001100110", "110"), -- i=324
      ("1001000001100110", "110"), -- i=325
      ("1010000001100110", "110"), -- i=326
      ("1011000001100110", "110"), -- i=327
      ("0101000001100000", "110"), -- i=328
      ("0100000001100000", "110"), -- i=329
      ("1000000001100111", "110"), -- i=330
      ("1001000001100111", "110"), -- i=331
      ("1010000001100111", "110"), -- i=332
      ("1011000001100111", "110"), -- i=333
      ("0101000001100000", "110"), -- i=334
      ("0100000001100000", "110"), -- i=335
      ("1000000001110000", "111"), -- i=336
      ("1001000001110000", "111"), -- i=337
      ("1010000001110000", "111"), -- i=338
      ("1011000001110000", "111"), -- i=339
      ("0101000001110000", "111"), -- i=340
      ("0100000001110000", "111"), -- i=341
      ("1000000001110001", "111"), -- i=342
      ("1001000001110001", "111"), -- i=343
      ("1010000001110001", "111"), -- i=344
      ("1011000001110001", "111"), -- i=345
      ("0101000001110000", "111"), -- i=346
      ("0100000001110000", "111"), -- i=347
      ("1000000001110010", "111"), -- i=348
      ("1001000001110010", "111"), -- i=349
      ("1010000001110010", "111"), -- i=350
      ("1011000001110010", "111"), -- i=351
      ("0101000001110000", "111"), -- i=352
      ("0100000001110000", "111"), -- i=353
      ("1000000001110011", "111"), -- i=354
      ("1001000001110011", "111"), -- i=355
      ("1010000001110011", "111"), -- i=356
      ("1011000001110011", "111"), -- i=357
      ("0101000001110000", "111"), -- i=358
      ("0100000001110000", "111"), -- i=359
      ("1000000001110100", "111"), -- i=360
      ("1001000001110100", "111"), -- i=361
      ("1010000001110100", "111"), -- i=362
      ("1011000001110100", "111"), -- i=363
      ("0101000001110000", "111"), -- i=364
      ("0100000001110000", "111"), -- i=365
      ("1000000001110101", "111"), -- i=366
      ("1001000001110101", "111"), -- i=367
      ("1010000001110101", "111"), -- i=368
      ("1011000001110101", "111"), -- i=369
      ("0101000001110000", "111"), -- i=370
      ("0100000001110000", "111"), -- i=371
      ("1000000001110110", "111"), -- i=372
      ("1001000001110110", "111"), -- i=373
      ("1010000001110110", "111"), -- i=374
      ("1011000001110110", "111"), -- i=375
      ("0101000001110000", "111"), -- i=376
      ("0100000001110000", "111"), -- i=377
      ("1000000001110111", "111"), -- i=378
      ("1001000001110111", "111"), -- i=379
      ("1010000001110111", "111"), -- i=380
      ("1011000001110111", "111"), -- i=381
      ("0101000001110000", "111"), -- i=382
      ("0100000001110000", "111"), -- i=383
      ("1000000100000000", "000"), -- i=384
      ("1001000100000000", "000"), -- i=385
      ("1010000100000000", "000"), -- i=386
      ("1011000100000000", "000"), -- i=387
      ("0101000100000000", "000"), -- i=388
      ("0100000100000000", "000"), -- i=389
      ("1000000100000001", "000"), -- i=390
      ("1001000100000001", "000"), -- i=391
      ("1010000100000001", "000"), -- i=392
      ("1011000100000001", "000"), -- i=393
      ("0101000100000000", "000"), -- i=394
      ("0100000100000000", "000"), -- i=395
      ("1000000100000010", "000"), -- i=396
      ("1001000100000010", "000"), -- i=397
      ("1010000100000010", "000"), -- i=398
      ("1011000100000010", "000"), -- i=399
      ("0101000100000000", "000"), -- i=400
      ("0100000100000000", "000"), -- i=401
      ("1000000100000011", "000"), -- i=402
      ("1001000100000011", "000"), -- i=403
      ("1010000100000011", "000"), -- i=404
      ("1011000100000011", "000"), -- i=405
      ("0101000100000000", "000"), -- i=406
      ("0100000100000000", "000"), -- i=407
      ("1000000100000100", "000"), -- i=408
      ("1001000100000100", "000"), -- i=409
      ("1010000100000100", "000"), -- i=410
      ("1011000100000100", "000"), -- i=411
      ("0101000100000000", "000"), -- i=412
      ("0100000100000000", "000"), -- i=413
      ("1000000100000101", "000"), -- i=414
      ("1001000100000101", "000"), -- i=415
      ("1010000100000101", "000"), -- i=416
      ("1011000100000101", "000"), -- i=417
      ("0101000100000000", "000"), -- i=418
      ("0100000100000000", "000"), -- i=419
      ("1000000100000110", "000"), -- i=420
      ("1001000100000110", "000"), -- i=421
      ("1010000100000110", "000"), -- i=422
      ("1011000100000110", "000"), -- i=423
      ("0101000100000000", "000"), -- i=424
      ("0100000100000000", "000"), -- i=425
      ("1000000100000111", "000"), -- i=426
      ("1001000100000111", "000"), -- i=427
      ("1010000100000111", "000"), -- i=428
      ("1011000100000111", "000"), -- i=429
      ("0101000100000000", "000"), -- i=430
      ("0100000100000000", "000"), -- i=431
      ("1000000100010000", "001"), -- i=432
      ("1001000100010000", "001"), -- i=433
      ("1010000100010000", "001"), -- i=434
      ("1011000100010000", "001"), -- i=435
      ("0101000100010000", "001"), -- i=436
      ("0100000100010000", "001"), -- i=437
      ("1000000100010001", "001"), -- i=438
      ("1001000100010001", "001"), -- i=439
      ("1010000100010001", "001"), -- i=440
      ("1011000100010001", "001"), -- i=441
      ("0101000100010000", "001"), -- i=442
      ("0100000100010000", "001"), -- i=443
      ("1000000100010010", "001"), -- i=444
      ("1001000100010010", "001"), -- i=445
      ("1010000100010010", "001"), -- i=446
      ("1011000100010010", "001"), -- i=447
      ("0101000100010000", "001"), -- i=448
      ("0100000100010000", "001"), -- i=449
      ("1000000100010011", "001"), -- i=450
      ("1001000100010011", "001"), -- i=451
      ("1010000100010011", "001"), -- i=452
      ("1011000100010011", "001"), -- i=453
      ("0101000100010000", "001"), -- i=454
      ("0100000100010000", "001"), -- i=455
      ("1000000100010100", "001"), -- i=456
      ("1001000100010100", "001"), -- i=457
      ("1010000100010100", "001"), -- i=458
      ("1011000100010100", "001"), -- i=459
      ("0101000100010000", "001"), -- i=460
      ("0100000100010000", "001"), -- i=461
      ("1000000100010101", "001"), -- i=462
      ("1001000100010101", "001"), -- i=463
      ("1010000100010101", "001"), -- i=464
      ("1011000100010101", "001"), -- i=465
      ("0101000100010000", "001"), -- i=466
      ("0100000100010000", "001"), -- i=467
      ("1000000100010110", "001"), -- i=468
      ("1001000100010110", "001"), -- i=469
      ("1010000100010110", "001"), -- i=470
      ("1011000100010110", "001"), -- i=471
      ("0101000100010000", "001"), -- i=472
      ("0100000100010000", "001"), -- i=473
      ("1000000100010111", "001"), -- i=474
      ("1001000100010111", "001"), -- i=475
      ("1010000100010111", "001"), -- i=476
      ("1011000100010111", "001"), -- i=477
      ("0101000100010000", "001"), -- i=478
      ("0100000100010000", "001"), -- i=479
      ("1000000100100000", "010"), -- i=480
      ("1001000100100000", "010"), -- i=481
      ("1010000100100000", "010"), -- i=482
      ("1011000100100000", "010"), -- i=483
      ("0101000100100000", "010"), -- i=484
      ("0100000100100000", "010"), -- i=485
      ("1000000100100001", "010"), -- i=486
      ("1001000100100001", "010"), -- i=487
      ("1010000100100001", "010"), -- i=488
      ("1011000100100001", "010"), -- i=489
      ("0101000100100000", "010"), -- i=490
      ("0100000100100000", "010"), -- i=491
      ("1000000100100010", "010"), -- i=492
      ("1001000100100010", "010"), -- i=493
      ("1010000100100010", "010"), -- i=494
      ("1011000100100010", "010"), -- i=495
      ("0101000100100000", "010"), -- i=496
      ("0100000100100000", "010"), -- i=497
      ("1000000100100011", "010"), -- i=498
      ("1001000100100011", "010"), -- i=499
      ("1010000100100011", "010"), -- i=500
      ("1011000100100011", "010"), -- i=501
      ("0101000100100000", "010"), -- i=502
      ("0100000100100000", "010"), -- i=503
      ("1000000100100100", "010"), -- i=504
      ("1001000100100100", "010"), -- i=505
      ("1010000100100100", "010"), -- i=506
      ("1011000100100100", "010"), -- i=507
      ("0101000100100000", "010"), -- i=508
      ("0100000100100000", "010"), -- i=509
      ("1000000100100101", "010"), -- i=510
      ("1001000100100101", "010"), -- i=511
      ("1010000100100101", "010"), -- i=512
      ("1011000100100101", "010"), -- i=513
      ("0101000100100000", "010"), -- i=514
      ("0100000100100000", "010"), -- i=515
      ("1000000100100110", "010"), -- i=516
      ("1001000100100110", "010"), -- i=517
      ("1010000100100110", "010"), -- i=518
      ("1011000100100110", "010"), -- i=519
      ("0101000100100000", "010"), -- i=520
      ("0100000100100000", "010"), -- i=521
      ("1000000100100111", "010"), -- i=522
      ("1001000100100111", "010"), -- i=523
      ("1010000100100111", "010"), -- i=524
      ("1011000100100111", "010"), -- i=525
      ("0101000100100000", "010"), -- i=526
      ("0100000100100000", "010"), -- i=527
      ("1000000100110000", "011"), -- i=528
      ("1001000100110000", "011"), -- i=529
      ("1010000100110000", "011"), -- i=530
      ("1011000100110000", "011"), -- i=531
      ("0101000100110000", "011"), -- i=532
      ("0100000100110000", "011"), -- i=533
      ("1000000100110001", "011"), -- i=534
      ("1001000100110001", "011"), -- i=535
      ("1010000100110001", "011"), -- i=536
      ("1011000100110001", "011"), -- i=537
      ("0101000100110000", "011"), -- i=538
      ("0100000100110000", "011"), -- i=539
      ("1000000100110010", "011"), -- i=540
      ("1001000100110010", "011"), -- i=541
      ("1010000100110010", "011"), -- i=542
      ("1011000100110010", "011"), -- i=543
      ("0101000100110000", "011"), -- i=544
      ("0100000100110000", "011"), -- i=545
      ("1000000100110011", "011"), -- i=546
      ("1001000100110011", "011"), -- i=547
      ("1010000100110011", "011"), -- i=548
      ("1011000100110011", "011"), -- i=549
      ("0101000100110000", "011"), -- i=550
      ("0100000100110000", "011"), -- i=551
      ("1000000100110100", "011"), -- i=552
      ("1001000100110100", "011"), -- i=553
      ("1010000100110100", "011"), -- i=554
      ("1011000100110100", "011"), -- i=555
      ("0101000100110000", "011"), -- i=556
      ("0100000100110000", "011"), -- i=557
      ("1000000100110101", "011"), -- i=558
      ("1001000100110101", "011"), -- i=559
      ("1010000100110101", "011"), -- i=560
      ("1011000100110101", "011"), -- i=561
      ("0101000100110000", "011"), -- i=562
      ("0100000100110000", "011"), -- i=563
      ("1000000100110110", "011"), -- i=564
      ("1001000100110110", "011"), -- i=565
      ("1010000100110110", "011"), -- i=566
      ("1011000100110110", "011"), -- i=567
      ("0101000100110000", "011"), -- i=568
      ("0100000100110000", "011"), -- i=569
      ("1000000100110111", "011"), -- i=570
      ("1001000100110111", "011"), -- i=571
      ("1010000100110111", "011"), -- i=572
      ("1011000100110111", "011"), -- i=573
      ("0101000100110000", "011"), -- i=574
      ("0100000100110000", "011"), -- i=575
      ("1000000101000000", "100"), -- i=576
      ("1001000101000000", "100"), -- i=577
      ("1010000101000000", "100"), -- i=578
      ("1011000101000000", "100"), -- i=579
      ("0101000101000000", "100"), -- i=580
      ("0100000101000000", "100"), -- i=581
      ("1000000101000001", "100"), -- i=582
      ("1001000101000001", "100"), -- i=583
      ("1010000101000001", "100"), -- i=584
      ("1011000101000001", "100"), -- i=585
      ("0101000101000000", "100"), -- i=586
      ("0100000101000000", "100"), -- i=587
      ("1000000101000010", "100"), -- i=588
      ("1001000101000010", "100"), -- i=589
      ("1010000101000010", "100"), -- i=590
      ("1011000101000010", "100"), -- i=591
      ("0101000101000000", "100"), -- i=592
      ("0100000101000000", "100"), -- i=593
      ("1000000101000011", "100"), -- i=594
      ("1001000101000011", "100"), -- i=595
      ("1010000101000011", "100"), -- i=596
      ("1011000101000011", "100"), -- i=597
      ("0101000101000000", "100"), -- i=598
      ("0100000101000000", "100"), -- i=599
      ("1000000101000100", "100"), -- i=600
      ("1001000101000100", "100"), -- i=601
      ("1010000101000100", "100"), -- i=602
      ("1011000101000100", "100"), -- i=603
      ("0101000101000000", "100"), -- i=604
      ("0100000101000000", "100"), -- i=605
      ("1000000101000101", "100"), -- i=606
      ("1001000101000101", "100"), -- i=607
      ("1010000101000101", "100"), -- i=608
      ("1011000101000101", "100"), -- i=609
      ("0101000101000000", "100"), -- i=610
      ("0100000101000000", "100"), -- i=611
      ("1000000101000110", "100"), -- i=612
      ("1001000101000110", "100"), -- i=613
      ("1010000101000110", "100"), -- i=614
      ("1011000101000110", "100"), -- i=615
      ("0101000101000000", "100"), -- i=616
      ("0100000101000000", "100"), -- i=617
      ("1000000101000111", "100"), -- i=618
      ("1001000101000111", "100"), -- i=619
      ("1010000101000111", "100"), -- i=620
      ("1011000101000111", "100"), -- i=621
      ("0101000101000000", "100"), -- i=622
      ("0100000101000000", "100"), -- i=623
      ("1000000101010000", "101"), -- i=624
      ("1001000101010000", "101"), -- i=625
      ("1010000101010000", "101"), -- i=626
      ("1011000101010000", "101"), -- i=627
      ("0101000101010000", "101"), -- i=628
      ("0100000101010000", "101"), -- i=629
      ("1000000101010001", "101"), -- i=630
      ("1001000101010001", "101"), -- i=631
      ("1010000101010001", "101"), -- i=632
      ("1011000101010001", "101"), -- i=633
      ("0101000101010000", "101"), -- i=634
      ("0100000101010000", "101"), -- i=635
      ("1000000101010010", "101"), -- i=636
      ("1001000101010010", "101"), -- i=637
      ("1010000101010010", "101"), -- i=638
      ("1011000101010010", "101"), -- i=639
      ("0101000101010000", "101"), -- i=640
      ("0100000101010000", "101"), -- i=641
      ("1000000101010011", "101"), -- i=642
      ("1001000101010011", "101"), -- i=643
      ("1010000101010011", "101"), -- i=644
      ("1011000101010011", "101"), -- i=645
      ("0101000101010000", "101"), -- i=646
      ("0100000101010000", "101"), -- i=647
      ("1000000101010100", "101"), -- i=648
      ("1001000101010100", "101"), -- i=649
      ("1010000101010100", "101"), -- i=650
      ("1011000101010100", "101"), -- i=651
      ("0101000101010000", "101"), -- i=652
      ("0100000101010000", "101"), -- i=653
      ("1000000101010101", "101"), -- i=654
      ("1001000101010101", "101"), -- i=655
      ("1010000101010101", "101"), -- i=656
      ("1011000101010101", "101"), -- i=657
      ("0101000101010000", "101"), -- i=658
      ("0100000101010000", "101"), -- i=659
      ("1000000101010110", "101"), -- i=660
      ("1001000101010110", "101"), -- i=661
      ("1010000101010110", "101"), -- i=662
      ("1011000101010110", "101"), -- i=663
      ("0101000101010000", "101"), -- i=664
      ("0100000101010000", "101"), -- i=665
      ("1000000101010111", "101"), -- i=666
      ("1001000101010111", "101"), -- i=667
      ("1010000101010111", "101"), -- i=668
      ("1011000101010111", "101"), -- i=669
      ("0101000101010000", "101"), -- i=670
      ("0100000101010000", "101"), -- i=671
      ("1000000101100000", "110"), -- i=672
      ("1001000101100000", "110"), -- i=673
      ("1010000101100000", "110"), -- i=674
      ("1011000101100000", "110"), -- i=675
      ("0101000101100000", "110"), -- i=676
      ("0100000101100000", "110"), -- i=677
      ("1000000101100001", "110"), -- i=678
      ("1001000101100001", "110"), -- i=679
      ("1010000101100001", "110"), -- i=680
      ("1011000101100001", "110"), -- i=681
      ("0101000101100000", "110"), -- i=682
      ("0100000101100000", "110"), -- i=683
      ("1000000101100010", "110"), -- i=684
      ("1001000101100010", "110"), -- i=685
      ("1010000101100010", "110"), -- i=686
      ("1011000101100010", "110"), -- i=687
      ("0101000101100000", "110"), -- i=688
      ("0100000101100000", "110"), -- i=689
      ("1000000101100011", "110"), -- i=690
      ("1001000101100011", "110"), -- i=691
      ("1010000101100011", "110"), -- i=692
      ("1011000101100011", "110"), -- i=693
      ("0101000101100000", "110"), -- i=694
      ("0100000101100000", "110"), -- i=695
      ("1000000101100100", "110"), -- i=696
      ("1001000101100100", "110"), -- i=697
      ("1010000101100100", "110"), -- i=698
      ("1011000101100100", "110"), -- i=699
      ("0101000101100000", "110"), -- i=700
      ("0100000101100000", "110"), -- i=701
      ("1000000101100101", "110"), -- i=702
      ("1001000101100101", "110"), -- i=703
      ("1010000101100101", "110"), -- i=704
      ("1011000101100101", "110"), -- i=705
      ("0101000101100000", "110"), -- i=706
      ("0100000101100000", "110"), -- i=707
      ("1000000101100110", "110"), -- i=708
      ("1001000101100110", "110"), -- i=709
      ("1010000101100110", "110"), -- i=710
      ("1011000101100110", "110"), -- i=711
      ("0101000101100000", "110"), -- i=712
      ("0100000101100000", "110"), -- i=713
      ("1000000101100111", "110"), -- i=714
      ("1001000101100111", "110"), -- i=715
      ("1010000101100111", "110"), -- i=716
      ("1011000101100111", "110"), -- i=717
      ("0101000101100000", "110"), -- i=718
      ("0100000101100000", "110"), -- i=719
      ("1000000101110000", "111"), -- i=720
      ("1001000101110000", "111"), -- i=721
      ("1010000101110000", "111"), -- i=722
      ("1011000101110000", "111"), -- i=723
      ("0101000101110000", "111"), -- i=724
      ("0100000101110000", "111"), -- i=725
      ("1000000101110001", "111"), -- i=726
      ("1001000101110001", "111"), -- i=727
      ("1010000101110001", "111"), -- i=728
      ("1011000101110001", "111"), -- i=729
      ("0101000101110000", "111"), -- i=730
      ("0100000101110000", "111"), -- i=731
      ("1000000101110010", "111"), -- i=732
      ("1001000101110010", "111"), -- i=733
      ("1010000101110010", "111"), -- i=734
      ("1011000101110010", "111"), -- i=735
      ("0101000101110000", "111"), -- i=736
      ("0100000101110000", "111"), -- i=737
      ("1000000101110011", "111"), -- i=738
      ("1001000101110011", "111"), -- i=739
      ("1010000101110011", "111"), -- i=740
      ("1011000101110011", "111"), -- i=741
      ("0101000101110000", "111"), -- i=742
      ("0100000101110000", "111"), -- i=743
      ("1000000101110100", "111"), -- i=744
      ("1001000101110100", "111"), -- i=745
      ("1010000101110100", "111"), -- i=746
      ("1011000101110100", "111"), -- i=747
      ("0101000101110000", "111"), -- i=748
      ("0100000101110000", "111"), -- i=749
      ("1000000101110101", "111"), -- i=750
      ("1001000101110101", "111"), -- i=751
      ("1010000101110101", "111"), -- i=752
      ("1011000101110101", "111"), -- i=753
      ("0101000101110000", "111"), -- i=754
      ("0100000101110000", "111"), -- i=755
      ("1000000101110110", "111"), -- i=756
      ("1001000101110110", "111"), -- i=757
      ("1010000101110110", "111"), -- i=758
      ("1011000101110110", "111"), -- i=759
      ("0101000101110000", "111"), -- i=760
      ("0100000101110000", "111"), -- i=761
      ("1000000101110111", "111"), -- i=762
      ("1001000101110111", "111"), -- i=763
      ("1010000101110111", "111"), -- i=764
      ("1011000101110111", "111"), -- i=765
      ("0101000101110000", "111"), -- i=766
      ("0100000101110000", "111"), -- i=767
      ("1000001000000000", "000"), -- i=768
      ("1001001000000000", "000"), -- i=769
      ("1010001000000000", "000"), -- i=770
      ("1011001000000000", "000"), -- i=771
      ("0101001000000000", "000"), -- i=772
      ("0100001000000000", "000"), -- i=773
      ("1000001000000001", "000"), -- i=774
      ("1001001000000001", "000"), -- i=775
      ("1010001000000001", "000"), -- i=776
      ("1011001000000001", "000"), -- i=777
      ("0101001000000000", "000"), -- i=778
      ("0100001000000000", "000"), -- i=779
      ("1000001000000010", "000"), -- i=780
      ("1001001000000010", "000"), -- i=781
      ("1010001000000010", "000"), -- i=782
      ("1011001000000010", "000"), -- i=783
      ("0101001000000000", "000"), -- i=784
      ("0100001000000000", "000"), -- i=785
      ("1000001000000011", "000"), -- i=786
      ("1001001000000011", "000"), -- i=787
      ("1010001000000011", "000"), -- i=788
      ("1011001000000011", "000"), -- i=789
      ("0101001000000000", "000"), -- i=790
      ("0100001000000000", "000"), -- i=791
      ("1000001000000100", "000"), -- i=792
      ("1001001000000100", "000"), -- i=793
      ("1010001000000100", "000"), -- i=794
      ("1011001000000100", "000"), -- i=795
      ("0101001000000000", "000"), -- i=796
      ("0100001000000000", "000"), -- i=797
      ("1000001000000101", "000"), -- i=798
      ("1001001000000101", "000"), -- i=799
      ("1010001000000101", "000"), -- i=800
      ("1011001000000101", "000"), -- i=801
      ("0101001000000000", "000"), -- i=802
      ("0100001000000000", "000"), -- i=803
      ("1000001000000110", "000"), -- i=804
      ("1001001000000110", "000"), -- i=805
      ("1010001000000110", "000"), -- i=806
      ("1011001000000110", "000"), -- i=807
      ("0101001000000000", "000"), -- i=808
      ("0100001000000000", "000"), -- i=809
      ("1000001000000111", "000"), -- i=810
      ("1001001000000111", "000"), -- i=811
      ("1010001000000111", "000"), -- i=812
      ("1011001000000111", "000"), -- i=813
      ("0101001000000000", "000"), -- i=814
      ("0100001000000000", "000"), -- i=815
      ("1000001000010000", "001"), -- i=816
      ("1001001000010000", "001"), -- i=817
      ("1010001000010000", "001"), -- i=818
      ("1011001000010000", "001"), -- i=819
      ("0101001000010000", "001"), -- i=820
      ("0100001000010000", "001"), -- i=821
      ("1000001000010001", "001"), -- i=822
      ("1001001000010001", "001"), -- i=823
      ("1010001000010001", "001"), -- i=824
      ("1011001000010001", "001"), -- i=825
      ("0101001000010000", "001"), -- i=826
      ("0100001000010000", "001"), -- i=827
      ("1000001000010010", "001"), -- i=828
      ("1001001000010010", "001"), -- i=829
      ("1010001000010010", "001"), -- i=830
      ("1011001000010010", "001"), -- i=831
      ("0101001000010000", "001"), -- i=832
      ("0100001000010000", "001"), -- i=833
      ("1000001000010011", "001"), -- i=834
      ("1001001000010011", "001"), -- i=835
      ("1010001000010011", "001"), -- i=836
      ("1011001000010011", "001"), -- i=837
      ("0101001000010000", "001"), -- i=838
      ("0100001000010000", "001"), -- i=839
      ("1000001000010100", "001"), -- i=840
      ("1001001000010100", "001"), -- i=841
      ("1010001000010100", "001"), -- i=842
      ("1011001000010100", "001"), -- i=843
      ("0101001000010000", "001"), -- i=844
      ("0100001000010000", "001"), -- i=845
      ("1000001000010101", "001"), -- i=846
      ("1001001000010101", "001"), -- i=847
      ("1010001000010101", "001"), -- i=848
      ("1011001000010101", "001"), -- i=849
      ("0101001000010000", "001"), -- i=850
      ("0100001000010000", "001"), -- i=851
      ("1000001000010110", "001"), -- i=852
      ("1001001000010110", "001"), -- i=853
      ("1010001000010110", "001"), -- i=854
      ("1011001000010110", "001"), -- i=855
      ("0101001000010000", "001"), -- i=856
      ("0100001000010000", "001"), -- i=857
      ("1000001000010111", "001"), -- i=858
      ("1001001000010111", "001"), -- i=859
      ("1010001000010111", "001"), -- i=860
      ("1011001000010111", "001"), -- i=861
      ("0101001000010000", "001"), -- i=862
      ("0100001000010000", "001"), -- i=863
      ("1000001000100000", "010"), -- i=864
      ("1001001000100000", "010"), -- i=865
      ("1010001000100000", "010"), -- i=866
      ("1011001000100000", "010"), -- i=867
      ("0101001000100000", "010"), -- i=868
      ("0100001000100000", "010"), -- i=869
      ("1000001000100001", "010"), -- i=870
      ("1001001000100001", "010"), -- i=871
      ("1010001000100001", "010"), -- i=872
      ("1011001000100001", "010"), -- i=873
      ("0101001000100000", "010"), -- i=874
      ("0100001000100000", "010"), -- i=875
      ("1000001000100010", "010"), -- i=876
      ("1001001000100010", "010"), -- i=877
      ("1010001000100010", "010"), -- i=878
      ("1011001000100010", "010"), -- i=879
      ("0101001000100000", "010"), -- i=880
      ("0100001000100000", "010"), -- i=881
      ("1000001000100011", "010"), -- i=882
      ("1001001000100011", "010"), -- i=883
      ("1010001000100011", "010"), -- i=884
      ("1011001000100011", "010"), -- i=885
      ("0101001000100000", "010"), -- i=886
      ("0100001000100000", "010"), -- i=887
      ("1000001000100100", "010"), -- i=888
      ("1001001000100100", "010"), -- i=889
      ("1010001000100100", "010"), -- i=890
      ("1011001000100100", "010"), -- i=891
      ("0101001000100000", "010"), -- i=892
      ("0100001000100000", "010"), -- i=893
      ("1000001000100101", "010"), -- i=894
      ("1001001000100101", "010"), -- i=895
      ("1010001000100101", "010"), -- i=896
      ("1011001000100101", "010"), -- i=897
      ("0101001000100000", "010"), -- i=898
      ("0100001000100000", "010"), -- i=899
      ("1000001000100110", "010"), -- i=900
      ("1001001000100110", "010"), -- i=901
      ("1010001000100110", "010"), -- i=902
      ("1011001000100110", "010"), -- i=903
      ("0101001000100000", "010"), -- i=904
      ("0100001000100000", "010"), -- i=905
      ("1000001000100111", "010"), -- i=906
      ("1001001000100111", "010"), -- i=907
      ("1010001000100111", "010"), -- i=908
      ("1011001000100111", "010"), -- i=909
      ("0101001000100000", "010"), -- i=910
      ("0100001000100000", "010"), -- i=911
      ("1000001000110000", "011"), -- i=912
      ("1001001000110000", "011"), -- i=913
      ("1010001000110000", "011"), -- i=914
      ("1011001000110000", "011"), -- i=915
      ("0101001000110000", "011"), -- i=916
      ("0100001000110000", "011"), -- i=917
      ("1000001000110001", "011"), -- i=918
      ("1001001000110001", "011"), -- i=919
      ("1010001000110001", "011"), -- i=920
      ("1011001000110001", "011"), -- i=921
      ("0101001000110000", "011"), -- i=922
      ("0100001000110000", "011"), -- i=923
      ("1000001000110010", "011"), -- i=924
      ("1001001000110010", "011"), -- i=925
      ("1010001000110010", "011"), -- i=926
      ("1011001000110010", "011"), -- i=927
      ("0101001000110000", "011"), -- i=928
      ("0100001000110000", "011"), -- i=929
      ("1000001000110011", "011"), -- i=930
      ("1001001000110011", "011"), -- i=931
      ("1010001000110011", "011"), -- i=932
      ("1011001000110011", "011"), -- i=933
      ("0101001000110000", "011"), -- i=934
      ("0100001000110000", "011"), -- i=935
      ("1000001000110100", "011"), -- i=936
      ("1001001000110100", "011"), -- i=937
      ("1010001000110100", "011"), -- i=938
      ("1011001000110100", "011"), -- i=939
      ("0101001000110000", "011"), -- i=940
      ("0100001000110000", "011"), -- i=941
      ("1000001000110101", "011"), -- i=942
      ("1001001000110101", "011"), -- i=943
      ("1010001000110101", "011"), -- i=944
      ("1011001000110101", "011"), -- i=945
      ("0101001000110000", "011"), -- i=946
      ("0100001000110000", "011"), -- i=947
      ("1000001000110110", "011"), -- i=948
      ("1001001000110110", "011"), -- i=949
      ("1010001000110110", "011"), -- i=950
      ("1011001000110110", "011"), -- i=951
      ("0101001000110000", "011"), -- i=952
      ("0100001000110000", "011"), -- i=953
      ("1000001000110111", "011"), -- i=954
      ("1001001000110111", "011"), -- i=955
      ("1010001000110111", "011"), -- i=956
      ("1011001000110111", "011"), -- i=957
      ("0101001000110000", "011"), -- i=958
      ("0100001000110000", "011"), -- i=959
      ("1000001001000000", "100"), -- i=960
      ("1001001001000000", "100"), -- i=961
      ("1010001001000000", "100"), -- i=962
      ("1011001001000000", "100"), -- i=963
      ("0101001001000000", "100"), -- i=964
      ("0100001001000000", "100"), -- i=965
      ("1000001001000001", "100"), -- i=966
      ("1001001001000001", "100"), -- i=967
      ("1010001001000001", "100"), -- i=968
      ("1011001001000001", "100"), -- i=969
      ("0101001001000000", "100"), -- i=970
      ("0100001001000000", "100"), -- i=971
      ("1000001001000010", "100"), -- i=972
      ("1001001001000010", "100"), -- i=973
      ("1010001001000010", "100"), -- i=974
      ("1011001001000010", "100"), -- i=975
      ("0101001001000000", "100"), -- i=976
      ("0100001001000000", "100"), -- i=977
      ("1000001001000011", "100"), -- i=978
      ("1001001001000011", "100"), -- i=979
      ("1010001001000011", "100"), -- i=980
      ("1011001001000011", "100"), -- i=981
      ("0101001001000000", "100"), -- i=982
      ("0100001001000000", "100"), -- i=983
      ("1000001001000100", "100"), -- i=984
      ("1001001001000100", "100"), -- i=985
      ("1010001001000100", "100"), -- i=986
      ("1011001001000100", "100"), -- i=987
      ("0101001001000000", "100"), -- i=988
      ("0100001001000000", "100"), -- i=989
      ("1000001001000101", "100"), -- i=990
      ("1001001001000101", "100"), -- i=991
      ("1010001001000101", "100"), -- i=992
      ("1011001001000101", "100"), -- i=993
      ("0101001001000000", "100"), -- i=994
      ("0100001001000000", "100"), -- i=995
      ("1000001001000110", "100"), -- i=996
      ("1001001001000110", "100"), -- i=997
      ("1010001001000110", "100"), -- i=998
      ("1011001001000110", "100"), -- i=999
      ("0101001001000000", "100"), -- i=1000
      ("0100001001000000", "100"), -- i=1001
      ("1000001001000111", "100"), -- i=1002
      ("1001001001000111", "100"), -- i=1003
      ("1010001001000111", "100"), -- i=1004
      ("1011001001000111", "100"), -- i=1005
      ("0101001001000000", "100"), -- i=1006
      ("0100001001000000", "100"), -- i=1007
      ("1000001001010000", "101"), -- i=1008
      ("1001001001010000", "101"), -- i=1009
      ("1010001001010000", "101"), -- i=1010
      ("1011001001010000", "101"), -- i=1011
      ("0101001001010000", "101"), -- i=1012
      ("0100001001010000", "101"), -- i=1013
      ("1000001001010001", "101"), -- i=1014
      ("1001001001010001", "101"), -- i=1015
      ("1010001001010001", "101"), -- i=1016
      ("1011001001010001", "101"), -- i=1017
      ("0101001001010000", "101"), -- i=1018
      ("0100001001010000", "101"), -- i=1019
      ("1000001001010010", "101"), -- i=1020
      ("1001001001010010", "101"), -- i=1021
      ("1010001001010010", "101"), -- i=1022
      ("1011001001010010", "101"), -- i=1023
      ("0101001001010000", "101"), -- i=1024
      ("0100001001010000", "101"), -- i=1025
      ("1000001001010011", "101"), -- i=1026
      ("1001001001010011", "101"), -- i=1027
      ("1010001001010011", "101"), -- i=1028
      ("1011001001010011", "101"), -- i=1029
      ("0101001001010000", "101"), -- i=1030
      ("0100001001010000", "101"), -- i=1031
      ("1000001001010100", "101"), -- i=1032
      ("1001001001010100", "101"), -- i=1033
      ("1010001001010100", "101"), -- i=1034
      ("1011001001010100", "101"), -- i=1035
      ("0101001001010000", "101"), -- i=1036
      ("0100001001010000", "101"), -- i=1037
      ("1000001001010101", "101"), -- i=1038
      ("1001001001010101", "101"), -- i=1039
      ("1010001001010101", "101"), -- i=1040
      ("1011001001010101", "101"), -- i=1041
      ("0101001001010000", "101"), -- i=1042
      ("0100001001010000", "101"), -- i=1043
      ("1000001001010110", "101"), -- i=1044
      ("1001001001010110", "101"), -- i=1045
      ("1010001001010110", "101"), -- i=1046
      ("1011001001010110", "101"), -- i=1047
      ("0101001001010000", "101"), -- i=1048
      ("0100001001010000", "101"), -- i=1049
      ("1000001001010111", "101"), -- i=1050
      ("1001001001010111", "101"), -- i=1051
      ("1010001001010111", "101"), -- i=1052
      ("1011001001010111", "101"), -- i=1053
      ("0101001001010000", "101"), -- i=1054
      ("0100001001010000", "101"), -- i=1055
      ("1000001001100000", "110"), -- i=1056
      ("1001001001100000", "110"), -- i=1057
      ("1010001001100000", "110"), -- i=1058
      ("1011001001100000", "110"), -- i=1059
      ("0101001001100000", "110"), -- i=1060
      ("0100001001100000", "110"), -- i=1061
      ("1000001001100001", "110"), -- i=1062
      ("1001001001100001", "110"), -- i=1063
      ("1010001001100001", "110"), -- i=1064
      ("1011001001100001", "110"), -- i=1065
      ("0101001001100000", "110"), -- i=1066
      ("0100001001100000", "110"), -- i=1067
      ("1000001001100010", "110"), -- i=1068
      ("1001001001100010", "110"), -- i=1069
      ("1010001001100010", "110"), -- i=1070
      ("1011001001100010", "110"), -- i=1071
      ("0101001001100000", "110"), -- i=1072
      ("0100001001100000", "110"), -- i=1073
      ("1000001001100011", "110"), -- i=1074
      ("1001001001100011", "110"), -- i=1075
      ("1010001001100011", "110"), -- i=1076
      ("1011001001100011", "110"), -- i=1077
      ("0101001001100000", "110"), -- i=1078
      ("0100001001100000", "110"), -- i=1079
      ("1000001001100100", "110"), -- i=1080
      ("1001001001100100", "110"), -- i=1081
      ("1010001001100100", "110"), -- i=1082
      ("1011001001100100", "110"), -- i=1083
      ("0101001001100000", "110"), -- i=1084
      ("0100001001100000", "110"), -- i=1085
      ("1000001001100101", "110"), -- i=1086
      ("1001001001100101", "110"), -- i=1087
      ("1010001001100101", "110"), -- i=1088
      ("1011001001100101", "110"), -- i=1089
      ("0101001001100000", "110"), -- i=1090
      ("0100001001100000", "110"), -- i=1091
      ("1000001001100110", "110"), -- i=1092
      ("1001001001100110", "110"), -- i=1093
      ("1010001001100110", "110"), -- i=1094
      ("1011001001100110", "110"), -- i=1095
      ("0101001001100000", "110"), -- i=1096
      ("0100001001100000", "110"), -- i=1097
      ("1000001001100111", "110"), -- i=1098
      ("1001001001100111", "110"), -- i=1099
      ("1010001001100111", "110"), -- i=1100
      ("1011001001100111", "110"), -- i=1101
      ("0101001001100000", "110"), -- i=1102
      ("0100001001100000", "110"), -- i=1103
      ("1000001001110000", "111"), -- i=1104
      ("1001001001110000", "111"), -- i=1105
      ("1010001001110000", "111"), -- i=1106
      ("1011001001110000", "111"), -- i=1107
      ("0101001001110000", "111"), -- i=1108
      ("0100001001110000", "111"), -- i=1109
      ("1000001001110001", "111"), -- i=1110
      ("1001001001110001", "111"), -- i=1111
      ("1010001001110001", "111"), -- i=1112
      ("1011001001110001", "111"), -- i=1113
      ("0101001001110000", "111"), -- i=1114
      ("0100001001110000", "111"), -- i=1115
      ("1000001001110010", "111"), -- i=1116
      ("1001001001110010", "111"), -- i=1117
      ("1010001001110010", "111"), -- i=1118
      ("1011001001110010", "111"), -- i=1119
      ("0101001001110000", "111"), -- i=1120
      ("0100001001110000", "111"), -- i=1121
      ("1000001001110011", "111"), -- i=1122
      ("1001001001110011", "111"), -- i=1123
      ("1010001001110011", "111"), -- i=1124
      ("1011001001110011", "111"), -- i=1125
      ("0101001001110000", "111"), -- i=1126
      ("0100001001110000", "111"), -- i=1127
      ("1000001001110100", "111"), -- i=1128
      ("1001001001110100", "111"), -- i=1129
      ("1010001001110100", "111"), -- i=1130
      ("1011001001110100", "111"), -- i=1131
      ("0101001001110000", "111"), -- i=1132
      ("0100001001110000", "111"), -- i=1133
      ("1000001001110101", "111"), -- i=1134
      ("1001001001110101", "111"), -- i=1135
      ("1010001001110101", "111"), -- i=1136
      ("1011001001110101", "111"), -- i=1137
      ("0101001001110000", "111"), -- i=1138
      ("0100001001110000", "111"), -- i=1139
      ("1000001001110110", "111"), -- i=1140
      ("1001001001110110", "111"), -- i=1141
      ("1010001001110110", "111"), -- i=1142
      ("1011001001110110", "111"), -- i=1143
      ("0101001001110000", "111"), -- i=1144
      ("0100001001110000", "111"), -- i=1145
      ("1000001001110111", "111"), -- i=1146
      ("1001001001110111", "111"), -- i=1147
      ("1010001001110111", "111"), -- i=1148
      ("1011001001110111", "111"), -- i=1149
      ("0101001001110000", "111"), -- i=1150
      ("0100001001110000", "111"), -- i=1151
      ("1000001100000000", "000"), -- i=1152
      ("1001001100000000", "000"), -- i=1153
      ("1010001100000000", "000"), -- i=1154
      ("1011001100000000", "000"), -- i=1155
      ("0101001100000000", "000"), -- i=1156
      ("0100001100000000", "000"), -- i=1157
      ("1000001100000001", "000"), -- i=1158
      ("1001001100000001", "000"), -- i=1159
      ("1010001100000001", "000"), -- i=1160
      ("1011001100000001", "000"), -- i=1161
      ("0101001100000000", "000"), -- i=1162
      ("0100001100000000", "000"), -- i=1163
      ("1000001100000010", "000"), -- i=1164
      ("1001001100000010", "000"), -- i=1165
      ("1010001100000010", "000"), -- i=1166
      ("1011001100000010", "000"), -- i=1167
      ("0101001100000000", "000"), -- i=1168
      ("0100001100000000", "000"), -- i=1169
      ("1000001100000011", "000"), -- i=1170
      ("1001001100000011", "000"), -- i=1171
      ("1010001100000011", "000"), -- i=1172
      ("1011001100000011", "000"), -- i=1173
      ("0101001100000000", "000"), -- i=1174
      ("0100001100000000", "000"), -- i=1175
      ("1000001100000100", "000"), -- i=1176
      ("1001001100000100", "000"), -- i=1177
      ("1010001100000100", "000"), -- i=1178
      ("1011001100000100", "000"), -- i=1179
      ("0101001100000000", "000"), -- i=1180
      ("0100001100000000", "000"), -- i=1181
      ("1000001100000101", "000"), -- i=1182
      ("1001001100000101", "000"), -- i=1183
      ("1010001100000101", "000"), -- i=1184
      ("1011001100000101", "000"), -- i=1185
      ("0101001100000000", "000"), -- i=1186
      ("0100001100000000", "000"), -- i=1187
      ("1000001100000110", "000"), -- i=1188
      ("1001001100000110", "000"), -- i=1189
      ("1010001100000110", "000"), -- i=1190
      ("1011001100000110", "000"), -- i=1191
      ("0101001100000000", "000"), -- i=1192
      ("0100001100000000", "000"), -- i=1193
      ("1000001100000111", "000"), -- i=1194
      ("1001001100000111", "000"), -- i=1195
      ("1010001100000111", "000"), -- i=1196
      ("1011001100000111", "000"), -- i=1197
      ("0101001100000000", "000"), -- i=1198
      ("0100001100000000", "000"), -- i=1199
      ("1000001100010000", "001"), -- i=1200
      ("1001001100010000", "001"), -- i=1201
      ("1010001100010000", "001"), -- i=1202
      ("1011001100010000", "001"), -- i=1203
      ("0101001100010000", "001"), -- i=1204
      ("0100001100010000", "001"), -- i=1205
      ("1000001100010001", "001"), -- i=1206
      ("1001001100010001", "001"), -- i=1207
      ("1010001100010001", "001"), -- i=1208
      ("1011001100010001", "001"), -- i=1209
      ("0101001100010000", "001"), -- i=1210
      ("0100001100010000", "001"), -- i=1211
      ("1000001100010010", "001"), -- i=1212
      ("1001001100010010", "001"), -- i=1213
      ("1010001100010010", "001"), -- i=1214
      ("1011001100010010", "001"), -- i=1215
      ("0101001100010000", "001"), -- i=1216
      ("0100001100010000", "001"), -- i=1217
      ("1000001100010011", "001"), -- i=1218
      ("1001001100010011", "001"), -- i=1219
      ("1010001100010011", "001"), -- i=1220
      ("1011001100010011", "001"), -- i=1221
      ("0101001100010000", "001"), -- i=1222
      ("0100001100010000", "001"), -- i=1223
      ("1000001100010100", "001"), -- i=1224
      ("1001001100010100", "001"), -- i=1225
      ("1010001100010100", "001"), -- i=1226
      ("1011001100010100", "001"), -- i=1227
      ("0101001100010000", "001"), -- i=1228
      ("0100001100010000", "001"), -- i=1229
      ("1000001100010101", "001"), -- i=1230
      ("1001001100010101", "001"), -- i=1231
      ("1010001100010101", "001"), -- i=1232
      ("1011001100010101", "001"), -- i=1233
      ("0101001100010000", "001"), -- i=1234
      ("0100001100010000", "001"), -- i=1235
      ("1000001100010110", "001"), -- i=1236
      ("1001001100010110", "001"), -- i=1237
      ("1010001100010110", "001"), -- i=1238
      ("1011001100010110", "001"), -- i=1239
      ("0101001100010000", "001"), -- i=1240
      ("0100001100010000", "001"), -- i=1241
      ("1000001100010111", "001"), -- i=1242
      ("1001001100010111", "001"), -- i=1243
      ("1010001100010111", "001"), -- i=1244
      ("1011001100010111", "001"), -- i=1245
      ("0101001100010000", "001"), -- i=1246
      ("0100001100010000", "001"), -- i=1247
      ("1000001100100000", "010"), -- i=1248
      ("1001001100100000", "010"), -- i=1249
      ("1010001100100000", "010"), -- i=1250
      ("1011001100100000", "010"), -- i=1251
      ("0101001100100000", "010"), -- i=1252
      ("0100001100100000", "010"), -- i=1253
      ("1000001100100001", "010"), -- i=1254
      ("1001001100100001", "010"), -- i=1255
      ("1010001100100001", "010"), -- i=1256
      ("1011001100100001", "010"), -- i=1257
      ("0101001100100000", "010"), -- i=1258
      ("0100001100100000", "010"), -- i=1259
      ("1000001100100010", "010"), -- i=1260
      ("1001001100100010", "010"), -- i=1261
      ("1010001100100010", "010"), -- i=1262
      ("1011001100100010", "010"), -- i=1263
      ("0101001100100000", "010"), -- i=1264
      ("0100001100100000", "010"), -- i=1265
      ("1000001100100011", "010"), -- i=1266
      ("1001001100100011", "010"), -- i=1267
      ("1010001100100011", "010"), -- i=1268
      ("1011001100100011", "010"), -- i=1269
      ("0101001100100000", "010"), -- i=1270
      ("0100001100100000", "010"), -- i=1271
      ("1000001100100100", "010"), -- i=1272
      ("1001001100100100", "010"), -- i=1273
      ("1010001100100100", "010"), -- i=1274
      ("1011001100100100", "010"), -- i=1275
      ("0101001100100000", "010"), -- i=1276
      ("0100001100100000", "010"), -- i=1277
      ("1000001100100101", "010"), -- i=1278
      ("1001001100100101", "010"), -- i=1279
      ("1010001100100101", "010"), -- i=1280
      ("1011001100100101", "010"), -- i=1281
      ("0101001100100000", "010"), -- i=1282
      ("0100001100100000", "010"), -- i=1283
      ("1000001100100110", "010"), -- i=1284
      ("1001001100100110", "010"), -- i=1285
      ("1010001100100110", "010"), -- i=1286
      ("1011001100100110", "010"), -- i=1287
      ("0101001100100000", "010"), -- i=1288
      ("0100001100100000", "010"), -- i=1289
      ("1000001100100111", "010"), -- i=1290
      ("1001001100100111", "010"), -- i=1291
      ("1010001100100111", "010"), -- i=1292
      ("1011001100100111", "010"), -- i=1293
      ("0101001100100000", "010"), -- i=1294
      ("0100001100100000", "010"), -- i=1295
      ("1000001100110000", "011"), -- i=1296
      ("1001001100110000", "011"), -- i=1297
      ("1010001100110000", "011"), -- i=1298
      ("1011001100110000", "011"), -- i=1299
      ("0101001100110000", "011"), -- i=1300
      ("0100001100110000", "011"), -- i=1301
      ("1000001100110001", "011"), -- i=1302
      ("1001001100110001", "011"), -- i=1303
      ("1010001100110001", "011"), -- i=1304
      ("1011001100110001", "011"), -- i=1305
      ("0101001100110000", "011"), -- i=1306
      ("0100001100110000", "011"), -- i=1307
      ("1000001100110010", "011"), -- i=1308
      ("1001001100110010", "011"), -- i=1309
      ("1010001100110010", "011"), -- i=1310
      ("1011001100110010", "011"), -- i=1311
      ("0101001100110000", "011"), -- i=1312
      ("0100001100110000", "011"), -- i=1313
      ("1000001100110011", "011"), -- i=1314
      ("1001001100110011", "011"), -- i=1315
      ("1010001100110011", "011"), -- i=1316
      ("1011001100110011", "011"), -- i=1317
      ("0101001100110000", "011"), -- i=1318
      ("0100001100110000", "011"), -- i=1319
      ("1000001100110100", "011"), -- i=1320
      ("1001001100110100", "011"), -- i=1321
      ("1010001100110100", "011"), -- i=1322
      ("1011001100110100", "011"), -- i=1323
      ("0101001100110000", "011"), -- i=1324
      ("0100001100110000", "011"), -- i=1325
      ("1000001100110101", "011"), -- i=1326
      ("1001001100110101", "011"), -- i=1327
      ("1010001100110101", "011"), -- i=1328
      ("1011001100110101", "011"), -- i=1329
      ("0101001100110000", "011"), -- i=1330
      ("0100001100110000", "011"), -- i=1331
      ("1000001100110110", "011"), -- i=1332
      ("1001001100110110", "011"), -- i=1333
      ("1010001100110110", "011"), -- i=1334
      ("1011001100110110", "011"), -- i=1335
      ("0101001100110000", "011"), -- i=1336
      ("0100001100110000", "011"), -- i=1337
      ("1000001100110111", "011"), -- i=1338
      ("1001001100110111", "011"), -- i=1339
      ("1010001100110111", "011"), -- i=1340
      ("1011001100110111", "011"), -- i=1341
      ("0101001100110000", "011"), -- i=1342
      ("0100001100110000", "011"), -- i=1343
      ("1000001101000000", "100"), -- i=1344
      ("1001001101000000", "100"), -- i=1345
      ("1010001101000000", "100"), -- i=1346
      ("1011001101000000", "100"), -- i=1347
      ("0101001101000000", "100"), -- i=1348
      ("0100001101000000", "100"), -- i=1349
      ("1000001101000001", "100"), -- i=1350
      ("1001001101000001", "100"), -- i=1351
      ("1010001101000001", "100"), -- i=1352
      ("1011001101000001", "100"), -- i=1353
      ("0101001101000000", "100"), -- i=1354
      ("0100001101000000", "100"), -- i=1355
      ("1000001101000010", "100"), -- i=1356
      ("1001001101000010", "100"), -- i=1357
      ("1010001101000010", "100"), -- i=1358
      ("1011001101000010", "100"), -- i=1359
      ("0101001101000000", "100"), -- i=1360
      ("0100001101000000", "100"), -- i=1361
      ("1000001101000011", "100"), -- i=1362
      ("1001001101000011", "100"), -- i=1363
      ("1010001101000011", "100"), -- i=1364
      ("1011001101000011", "100"), -- i=1365
      ("0101001101000000", "100"), -- i=1366
      ("0100001101000000", "100"), -- i=1367
      ("1000001101000100", "100"), -- i=1368
      ("1001001101000100", "100"), -- i=1369
      ("1010001101000100", "100"), -- i=1370
      ("1011001101000100", "100"), -- i=1371
      ("0101001101000000", "100"), -- i=1372
      ("0100001101000000", "100"), -- i=1373
      ("1000001101000101", "100"), -- i=1374
      ("1001001101000101", "100"), -- i=1375
      ("1010001101000101", "100"), -- i=1376
      ("1011001101000101", "100"), -- i=1377
      ("0101001101000000", "100"), -- i=1378
      ("0100001101000000", "100"), -- i=1379
      ("1000001101000110", "100"), -- i=1380
      ("1001001101000110", "100"), -- i=1381
      ("1010001101000110", "100"), -- i=1382
      ("1011001101000110", "100"), -- i=1383
      ("0101001101000000", "100"), -- i=1384
      ("0100001101000000", "100"), -- i=1385
      ("1000001101000111", "100"), -- i=1386
      ("1001001101000111", "100"), -- i=1387
      ("1010001101000111", "100"), -- i=1388
      ("1011001101000111", "100"), -- i=1389
      ("0101001101000000", "100"), -- i=1390
      ("0100001101000000", "100"), -- i=1391
      ("1000001101010000", "101"), -- i=1392
      ("1001001101010000", "101"), -- i=1393
      ("1010001101010000", "101"), -- i=1394
      ("1011001101010000", "101"), -- i=1395
      ("0101001101010000", "101"), -- i=1396
      ("0100001101010000", "101"), -- i=1397
      ("1000001101010001", "101"), -- i=1398
      ("1001001101010001", "101"), -- i=1399
      ("1010001101010001", "101"), -- i=1400
      ("1011001101010001", "101"), -- i=1401
      ("0101001101010000", "101"), -- i=1402
      ("0100001101010000", "101"), -- i=1403
      ("1000001101010010", "101"), -- i=1404
      ("1001001101010010", "101"), -- i=1405
      ("1010001101010010", "101"), -- i=1406
      ("1011001101010010", "101"), -- i=1407
      ("0101001101010000", "101"), -- i=1408
      ("0100001101010000", "101"), -- i=1409
      ("1000001101010011", "101"), -- i=1410
      ("1001001101010011", "101"), -- i=1411
      ("1010001101010011", "101"), -- i=1412
      ("1011001101010011", "101"), -- i=1413
      ("0101001101010000", "101"), -- i=1414
      ("0100001101010000", "101"), -- i=1415
      ("1000001101010100", "101"), -- i=1416
      ("1001001101010100", "101"), -- i=1417
      ("1010001101010100", "101"), -- i=1418
      ("1011001101010100", "101"), -- i=1419
      ("0101001101010000", "101"), -- i=1420
      ("0100001101010000", "101"), -- i=1421
      ("1000001101010101", "101"), -- i=1422
      ("1001001101010101", "101"), -- i=1423
      ("1010001101010101", "101"), -- i=1424
      ("1011001101010101", "101"), -- i=1425
      ("0101001101010000", "101"), -- i=1426
      ("0100001101010000", "101"), -- i=1427
      ("1000001101010110", "101"), -- i=1428
      ("1001001101010110", "101"), -- i=1429
      ("1010001101010110", "101"), -- i=1430
      ("1011001101010110", "101"), -- i=1431
      ("0101001101010000", "101"), -- i=1432
      ("0100001101010000", "101"), -- i=1433
      ("1000001101010111", "101"), -- i=1434
      ("1001001101010111", "101"), -- i=1435
      ("1010001101010111", "101"), -- i=1436
      ("1011001101010111", "101"), -- i=1437
      ("0101001101010000", "101"), -- i=1438
      ("0100001101010000", "101"), -- i=1439
      ("1000001101100000", "110"), -- i=1440
      ("1001001101100000", "110"), -- i=1441
      ("1010001101100000", "110"), -- i=1442
      ("1011001101100000", "110"), -- i=1443
      ("0101001101100000", "110"), -- i=1444
      ("0100001101100000", "110"), -- i=1445
      ("1000001101100001", "110"), -- i=1446
      ("1001001101100001", "110"), -- i=1447
      ("1010001101100001", "110"), -- i=1448
      ("1011001101100001", "110"), -- i=1449
      ("0101001101100000", "110"), -- i=1450
      ("0100001101100000", "110"), -- i=1451
      ("1000001101100010", "110"), -- i=1452
      ("1001001101100010", "110"), -- i=1453
      ("1010001101100010", "110"), -- i=1454
      ("1011001101100010", "110"), -- i=1455
      ("0101001101100000", "110"), -- i=1456
      ("0100001101100000", "110"), -- i=1457
      ("1000001101100011", "110"), -- i=1458
      ("1001001101100011", "110"), -- i=1459
      ("1010001101100011", "110"), -- i=1460
      ("1011001101100011", "110"), -- i=1461
      ("0101001101100000", "110"), -- i=1462
      ("0100001101100000", "110"), -- i=1463
      ("1000001101100100", "110"), -- i=1464
      ("1001001101100100", "110"), -- i=1465
      ("1010001101100100", "110"), -- i=1466
      ("1011001101100100", "110"), -- i=1467
      ("0101001101100000", "110"), -- i=1468
      ("0100001101100000", "110"), -- i=1469
      ("1000001101100101", "110"), -- i=1470
      ("1001001101100101", "110"), -- i=1471
      ("1010001101100101", "110"), -- i=1472
      ("1011001101100101", "110"), -- i=1473
      ("0101001101100000", "110"), -- i=1474
      ("0100001101100000", "110"), -- i=1475
      ("1000001101100110", "110"), -- i=1476
      ("1001001101100110", "110"), -- i=1477
      ("1010001101100110", "110"), -- i=1478
      ("1011001101100110", "110"), -- i=1479
      ("0101001101100000", "110"), -- i=1480
      ("0100001101100000", "110"), -- i=1481
      ("1000001101100111", "110"), -- i=1482
      ("1001001101100111", "110"), -- i=1483
      ("1010001101100111", "110"), -- i=1484
      ("1011001101100111", "110"), -- i=1485
      ("0101001101100000", "110"), -- i=1486
      ("0100001101100000", "110"), -- i=1487
      ("1000001101110000", "111"), -- i=1488
      ("1001001101110000", "111"), -- i=1489
      ("1010001101110000", "111"), -- i=1490
      ("1011001101110000", "111"), -- i=1491
      ("0101001101110000", "111"), -- i=1492
      ("0100001101110000", "111"), -- i=1493
      ("1000001101110001", "111"), -- i=1494
      ("1001001101110001", "111"), -- i=1495
      ("1010001101110001", "111"), -- i=1496
      ("1011001101110001", "111"), -- i=1497
      ("0101001101110000", "111"), -- i=1498
      ("0100001101110000", "111"), -- i=1499
      ("1000001101110010", "111"), -- i=1500
      ("1001001101110010", "111"), -- i=1501
      ("1010001101110010", "111"), -- i=1502
      ("1011001101110010", "111"), -- i=1503
      ("0101001101110000", "111"), -- i=1504
      ("0100001101110000", "111"), -- i=1505
      ("1000001101110011", "111"), -- i=1506
      ("1001001101110011", "111"), -- i=1507
      ("1010001101110011", "111"), -- i=1508
      ("1011001101110011", "111"), -- i=1509
      ("0101001101110000", "111"), -- i=1510
      ("0100001101110000", "111"), -- i=1511
      ("1000001101110100", "111"), -- i=1512
      ("1001001101110100", "111"), -- i=1513
      ("1010001101110100", "111"), -- i=1514
      ("1011001101110100", "111"), -- i=1515
      ("0101001101110000", "111"), -- i=1516
      ("0100001101110000", "111"), -- i=1517
      ("1000001101110101", "111"), -- i=1518
      ("1001001101110101", "111"), -- i=1519
      ("1010001101110101", "111"), -- i=1520
      ("1011001101110101", "111"), -- i=1521
      ("0101001101110000", "111"), -- i=1522
      ("0100001101110000", "111"), -- i=1523
      ("1000001101110110", "111"), -- i=1524
      ("1001001101110110", "111"), -- i=1525
      ("1010001101110110", "111"), -- i=1526
      ("1011001101110110", "111"), -- i=1527
      ("0101001101110000", "111"), -- i=1528
      ("0100001101110000", "111"), -- i=1529
      ("1000001101110111", "111"), -- i=1530
      ("1001001101110111", "111"), -- i=1531
      ("1010001101110111", "111"), -- i=1532
      ("1011001101110111", "111"), -- i=1533
      ("0101001101110000", "111"), -- i=1534
      ("0100001101110000", "111"), -- i=1535
      ("1000010000000000", "000"), -- i=1536
      ("1001010000000000", "000"), -- i=1537
      ("1010010000000000", "000"), -- i=1538
      ("1011010000000000", "000"), -- i=1539
      ("0101010000000000", "000"), -- i=1540
      ("0100010000000000", "000"), -- i=1541
      ("1000010000000001", "000"), -- i=1542
      ("1001010000000001", "000"), -- i=1543
      ("1010010000000001", "000"), -- i=1544
      ("1011010000000001", "000"), -- i=1545
      ("0101010000000000", "000"), -- i=1546
      ("0100010000000000", "000"), -- i=1547
      ("1000010000000010", "000"), -- i=1548
      ("1001010000000010", "000"), -- i=1549
      ("1010010000000010", "000"), -- i=1550
      ("1011010000000010", "000"), -- i=1551
      ("0101010000000000", "000"), -- i=1552
      ("0100010000000000", "000"), -- i=1553
      ("1000010000000011", "000"), -- i=1554
      ("1001010000000011", "000"), -- i=1555
      ("1010010000000011", "000"), -- i=1556
      ("1011010000000011", "000"), -- i=1557
      ("0101010000000000", "000"), -- i=1558
      ("0100010000000000", "000"), -- i=1559
      ("1000010000000100", "000"), -- i=1560
      ("1001010000000100", "000"), -- i=1561
      ("1010010000000100", "000"), -- i=1562
      ("1011010000000100", "000"), -- i=1563
      ("0101010000000000", "000"), -- i=1564
      ("0100010000000000", "000"), -- i=1565
      ("1000010000000101", "000"), -- i=1566
      ("1001010000000101", "000"), -- i=1567
      ("1010010000000101", "000"), -- i=1568
      ("1011010000000101", "000"), -- i=1569
      ("0101010000000000", "000"), -- i=1570
      ("0100010000000000", "000"), -- i=1571
      ("1000010000000110", "000"), -- i=1572
      ("1001010000000110", "000"), -- i=1573
      ("1010010000000110", "000"), -- i=1574
      ("1011010000000110", "000"), -- i=1575
      ("0101010000000000", "000"), -- i=1576
      ("0100010000000000", "000"), -- i=1577
      ("1000010000000111", "000"), -- i=1578
      ("1001010000000111", "000"), -- i=1579
      ("1010010000000111", "000"), -- i=1580
      ("1011010000000111", "000"), -- i=1581
      ("0101010000000000", "000"), -- i=1582
      ("0100010000000000", "000"), -- i=1583
      ("1000010000010000", "001"), -- i=1584
      ("1001010000010000", "001"), -- i=1585
      ("1010010000010000", "001"), -- i=1586
      ("1011010000010000", "001"), -- i=1587
      ("0101010000010000", "001"), -- i=1588
      ("0100010000010000", "001"), -- i=1589
      ("1000010000010001", "001"), -- i=1590
      ("1001010000010001", "001"), -- i=1591
      ("1010010000010001", "001"), -- i=1592
      ("1011010000010001", "001"), -- i=1593
      ("0101010000010000", "001"), -- i=1594
      ("0100010000010000", "001"), -- i=1595
      ("1000010000010010", "001"), -- i=1596
      ("1001010000010010", "001"), -- i=1597
      ("1010010000010010", "001"), -- i=1598
      ("1011010000010010", "001"), -- i=1599
      ("0101010000010000", "001"), -- i=1600
      ("0100010000010000", "001"), -- i=1601
      ("1000010000010011", "001"), -- i=1602
      ("1001010000010011", "001"), -- i=1603
      ("1010010000010011", "001"), -- i=1604
      ("1011010000010011", "001"), -- i=1605
      ("0101010000010000", "001"), -- i=1606
      ("0100010000010000", "001"), -- i=1607
      ("1000010000010100", "001"), -- i=1608
      ("1001010000010100", "001"), -- i=1609
      ("1010010000010100", "001"), -- i=1610
      ("1011010000010100", "001"), -- i=1611
      ("0101010000010000", "001"), -- i=1612
      ("0100010000010000", "001"), -- i=1613
      ("1000010000010101", "001"), -- i=1614
      ("1001010000010101", "001"), -- i=1615
      ("1010010000010101", "001"), -- i=1616
      ("1011010000010101", "001"), -- i=1617
      ("0101010000010000", "001"), -- i=1618
      ("0100010000010000", "001"), -- i=1619
      ("1000010000010110", "001"), -- i=1620
      ("1001010000010110", "001"), -- i=1621
      ("1010010000010110", "001"), -- i=1622
      ("1011010000010110", "001"), -- i=1623
      ("0101010000010000", "001"), -- i=1624
      ("0100010000010000", "001"), -- i=1625
      ("1000010000010111", "001"), -- i=1626
      ("1001010000010111", "001"), -- i=1627
      ("1010010000010111", "001"), -- i=1628
      ("1011010000010111", "001"), -- i=1629
      ("0101010000010000", "001"), -- i=1630
      ("0100010000010000", "001"), -- i=1631
      ("1000010000100000", "010"), -- i=1632
      ("1001010000100000", "010"), -- i=1633
      ("1010010000100000", "010"), -- i=1634
      ("1011010000100000", "010"), -- i=1635
      ("0101010000100000", "010"), -- i=1636
      ("0100010000100000", "010"), -- i=1637
      ("1000010000100001", "010"), -- i=1638
      ("1001010000100001", "010"), -- i=1639
      ("1010010000100001", "010"), -- i=1640
      ("1011010000100001", "010"), -- i=1641
      ("0101010000100000", "010"), -- i=1642
      ("0100010000100000", "010"), -- i=1643
      ("1000010000100010", "010"), -- i=1644
      ("1001010000100010", "010"), -- i=1645
      ("1010010000100010", "010"), -- i=1646
      ("1011010000100010", "010"), -- i=1647
      ("0101010000100000", "010"), -- i=1648
      ("0100010000100000", "010"), -- i=1649
      ("1000010000100011", "010"), -- i=1650
      ("1001010000100011", "010"), -- i=1651
      ("1010010000100011", "010"), -- i=1652
      ("1011010000100011", "010"), -- i=1653
      ("0101010000100000", "010"), -- i=1654
      ("0100010000100000", "010"), -- i=1655
      ("1000010000100100", "010"), -- i=1656
      ("1001010000100100", "010"), -- i=1657
      ("1010010000100100", "010"), -- i=1658
      ("1011010000100100", "010"), -- i=1659
      ("0101010000100000", "010"), -- i=1660
      ("0100010000100000", "010"), -- i=1661
      ("1000010000100101", "010"), -- i=1662
      ("1001010000100101", "010"), -- i=1663
      ("1010010000100101", "010"), -- i=1664
      ("1011010000100101", "010"), -- i=1665
      ("0101010000100000", "010"), -- i=1666
      ("0100010000100000", "010"), -- i=1667
      ("1000010000100110", "010"), -- i=1668
      ("1001010000100110", "010"), -- i=1669
      ("1010010000100110", "010"), -- i=1670
      ("1011010000100110", "010"), -- i=1671
      ("0101010000100000", "010"), -- i=1672
      ("0100010000100000", "010"), -- i=1673
      ("1000010000100111", "010"), -- i=1674
      ("1001010000100111", "010"), -- i=1675
      ("1010010000100111", "010"), -- i=1676
      ("1011010000100111", "010"), -- i=1677
      ("0101010000100000", "010"), -- i=1678
      ("0100010000100000", "010"), -- i=1679
      ("1000010000110000", "011"), -- i=1680
      ("1001010000110000", "011"), -- i=1681
      ("1010010000110000", "011"), -- i=1682
      ("1011010000110000", "011"), -- i=1683
      ("0101010000110000", "011"), -- i=1684
      ("0100010000110000", "011"), -- i=1685
      ("1000010000110001", "011"), -- i=1686
      ("1001010000110001", "011"), -- i=1687
      ("1010010000110001", "011"), -- i=1688
      ("1011010000110001", "011"), -- i=1689
      ("0101010000110000", "011"), -- i=1690
      ("0100010000110000", "011"), -- i=1691
      ("1000010000110010", "011"), -- i=1692
      ("1001010000110010", "011"), -- i=1693
      ("1010010000110010", "011"), -- i=1694
      ("1011010000110010", "011"), -- i=1695
      ("0101010000110000", "011"), -- i=1696
      ("0100010000110000", "011"), -- i=1697
      ("1000010000110011", "011"), -- i=1698
      ("1001010000110011", "011"), -- i=1699
      ("1010010000110011", "011"), -- i=1700
      ("1011010000110011", "011"), -- i=1701
      ("0101010000110000", "011"), -- i=1702
      ("0100010000110000", "011"), -- i=1703
      ("1000010000110100", "011"), -- i=1704
      ("1001010000110100", "011"), -- i=1705
      ("1010010000110100", "011"), -- i=1706
      ("1011010000110100", "011"), -- i=1707
      ("0101010000110000", "011"), -- i=1708
      ("0100010000110000", "011"), -- i=1709
      ("1000010000110101", "011"), -- i=1710
      ("1001010000110101", "011"), -- i=1711
      ("1010010000110101", "011"), -- i=1712
      ("1011010000110101", "011"), -- i=1713
      ("0101010000110000", "011"), -- i=1714
      ("0100010000110000", "011"), -- i=1715
      ("1000010000110110", "011"), -- i=1716
      ("1001010000110110", "011"), -- i=1717
      ("1010010000110110", "011"), -- i=1718
      ("1011010000110110", "011"), -- i=1719
      ("0101010000110000", "011"), -- i=1720
      ("0100010000110000", "011"), -- i=1721
      ("1000010000110111", "011"), -- i=1722
      ("1001010000110111", "011"), -- i=1723
      ("1010010000110111", "011"), -- i=1724
      ("1011010000110111", "011"), -- i=1725
      ("0101010000110000", "011"), -- i=1726
      ("0100010000110000", "011"), -- i=1727
      ("1000010001000000", "100"), -- i=1728
      ("1001010001000000", "100"), -- i=1729
      ("1010010001000000", "100"), -- i=1730
      ("1011010001000000", "100"), -- i=1731
      ("0101010001000000", "100"), -- i=1732
      ("0100010001000000", "100"), -- i=1733
      ("1000010001000001", "100"), -- i=1734
      ("1001010001000001", "100"), -- i=1735
      ("1010010001000001", "100"), -- i=1736
      ("1011010001000001", "100"), -- i=1737
      ("0101010001000000", "100"), -- i=1738
      ("0100010001000000", "100"), -- i=1739
      ("1000010001000010", "100"), -- i=1740
      ("1001010001000010", "100"), -- i=1741
      ("1010010001000010", "100"), -- i=1742
      ("1011010001000010", "100"), -- i=1743
      ("0101010001000000", "100"), -- i=1744
      ("0100010001000000", "100"), -- i=1745
      ("1000010001000011", "100"), -- i=1746
      ("1001010001000011", "100"), -- i=1747
      ("1010010001000011", "100"), -- i=1748
      ("1011010001000011", "100"), -- i=1749
      ("0101010001000000", "100"), -- i=1750
      ("0100010001000000", "100"), -- i=1751
      ("1000010001000100", "100"), -- i=1752
      ("1001010001000100", "100"), -- i=1753
      ("1010010001000100", "100"), -- i=1754
      ("1011010001000100", "100"), -- i=1755
      ("0101010001000000", "100"), -- i=1756
      ("0100010001000000", "100"), -- i=1757
      ("1000010001000101", "100"), -- i=1758
      ("1001010001000101", "100"), -- i=1759
      ("1010010001000101", "100"), -- i=1760
      ("1011010001000101", "100"), -- i=1761
      ("0101010001000000", "100"), -- i=1762
      ("0100010001000000", "100"), -- i=1763
      ("1000010001000110", "100"), -- i=1764
      ("1001010001000110", "100"), -- i=1765
      ("1010010001000110", "100"), -- i=1766
      ("1011010001000110", "100"), -- i=1767
      ("0101010001000000", "100"), -- i=1768
      ("0100010001000000", "100"), -- i=1769
      ("1000010001000111", "100"), -- i=1770
      ("1001010001000111", "100"), -- i=1771
      ("1010010001000111", "100"), -- i=1772
      ("1011010001000111", "100"), -- i=1773
      ("0101010001000000", "100"), -- i=1774
      ("0100010001000000", "100"), -- i=1775
      ("1000010001010000", "101"), -- i=1776
      ("1001010001010000", "101"), -- i=1777
      ("1010010001010000", "101"), -- i=1778
      ("1011010001010000", "101"), -- i=1779
      ("0101010001010000", "101"), -- i=1780
      ("0100010001010000", "101"), -- i=1781
      ("1000010001010001", "101"), -- i=1782
      ("1001010001010001", "101"), -- i=1783
      ("1010010001010001", "101"), -- i=1784
      ("1011010001010001", "101"), -- i=1785
      ("0101010001010000", "101"), -- i=1786
      ("0100010001010000", "101"), -- i=1787
      ("1000010001010010", "101"), -- i=1788
      ("1001010001010010", "101"), -- i=1789
      ("1010010001010010", "101"), -- i=1790
      ("1011010001010010", "101"), -- i=1791
      ("0101010001010000", "101"), -- i=1792
      ("0100010001010000", "101"), -- i=1793
      ("1000010001010011", "101"), -- i=1794
      ("1001010001010011", "101"), -- i=1795
      ("1010010001010011", "101"), -- i=1796
      ("1011010001010011", "101"), -- i=1797
      ("0101010001010000", "101"), -- i=1798
      ("0100010001010000", "101"), -- i=1799
      ("1000010001010100", "101"), -- i=1800
      ("1001010001010100", "101"), -- i=1801
      ("1010010001010100", "101"), -- i=1802
      ("1011010001010100", "101"), -- i=1803
      ("0101010001010000", "101"), -- i=1804
      ("0100010001010000", "101"), -- i=1805
      ("1000010001010101", "101"), -- i=1806
      ("1001010001010101", "101"), -- i=1807
      ("1010010001010101", "101"), -- i=1808
      ("1011010001010101", "101"), -- i=1809
      ("0101010001010000", "101"), -- i=1810
      ("0100010001010000", "101"), -- i=1811
      ("1000010001010110", "101"), -- i=1812
      ("1001010001010110", "101"), -- i=1813
      ("1010010001010110", "101"), -- i=1814
      ("1011010001010110", "101"), -- i=1815
      ("0101010001010000", "101"), -- i=1816
      ("0100010001010000", "101"), -- i=1817
      ("1000010001010111", "101"), -- i=1818
      ("1001010001010111", "101"), -- i=1819
      ("1010010001010111", "101"), -- i=1820
      ("1011010001010111", "101"), -- i=1821
      ("0101010001010000", "101"), -- i=1822
      ("0100010001010000", "101"), -- i=1823
      ("1000010001100000", "110"), -- i=1824
      ("1001010001100000", "110"), -- i=1825
      ("1010010001100000", "110"), -- i=1826
      ("1011010001100000", "110"), -- i=1827
      ("0101010001100000", "110"), -- i=1828
      ("0100010001100000", "110"), -- i=1829
      ("1000010001100001", "110"), -- i=1830
      ("1001010001100001", "110"), -- i=1831
      ("1010010001100001", "110"), -- i=1832
      ("1011010001100001", "110"), -- i=1833
      ("0101010001100000", "110"), -- i=1834
      ("0100010001100000", "110"), -- i=1835
      ("1000010001100010", "110"), -- i=1836
      ("1001010001100010", "110"), -- i=1837
      ("1010010001100010", "110"), -- i=1838
      ("1011010001100010", "110"), -- i=1839
      ("0101010001100000", "110"), -- i=1840
      ("0100010001100000", "110"), -- i=1841
      ("1000010001100011", "110"), -- i=1842
      ("1001010001100011", "110"), -- i=1843
      ("1010010001100011", "110"), -- i=1844
      ("1011010001100011", "110"), -- i=1845
      ("0101010001100000", "110"), -- i=1846
      ("0100010001100000", "110"), -- i=1847
      ("1000010001100100", "110"), -- i=1848
      ("1001010001100100", "110"), -- i=1849
      ("1010010001100100", "110"), -- i=1850
      ("1011010001100100", "110"), -- i=1851
      ("0101010001100000", "110"), -- i=1852
      ("0100010001100000", "110"), -- i=1853
      ("1000010001100101", "110"), -- i=1854
      ("1001010001100101", "110"), -- i=1855
      ("1010010001100101", "110"), -- i=1856
      ("1011010001100101", "110"), -- i=1857
      ("0101010001100000", "110"), -- i=1858
      ("0100010001100000", "110"), -- i=1859
      ("1000010001100110", "110"), -- i=1860
      ("1001010001100110", "110"), -- i=1861
      ("1010010001100110", "110"), -- i=1862
      ("1011010001100110", "110"), -- i=1863
      ("0101010001100000", "110"), -- i=1864
      ("0100010001100000", "110"), -- i=1865
      ("1000010001100111", "110"), -- i=1866
      ("1001010001100111", "110"), -- i=1867
      ("1010010001100111", "110"), -- i=1868
      ("1011010001100111", "110"), -- i=1869
      ("0101010001100000", "110"), -- i=1870
      ("0100010001100000", "110"), -- i=1871
      ("1000010001110000", "111"), -- i=1872
      ("1001010001110000", "111"), -- i=1873
      ("1010010001110000", "111"), -- i=1874
      ("1011010001110000", "111"), -- i=1875
      ("0101010001110000", "111"), -- i=1876
      ("0100010001110000", "111"), -- i=1877
      ("1000010001110001", "111"), -- i=1878
      ("1001010001110001", "111"), -- i=1879
      ("1010010001110001", "111"), -- i=1880
      ("1011010001110001", "111"), -- i=1881
      ("0101010001110000", "111"), -- i=1882
      ("0100010001110000", "111"), -- i=1883
      ("1000010001110010", "111"), -- i=1884
      ("1001010001110010", "111"), -- i=1885
      ("1010010001110010", "111"), -- i=1886
      ("1011010001110010", "111"), -- i=1887
      ("0101010001110000", "111"), -- i=1888
      ("0100010001110000", "111"), -- i=1889
      ("1000010001110011", "111"), -- i=1890
      ("1001010001110011", "111"), -- i=1891
      ("1010010001110011", "111"), -- i=1892
      ("1011010001110011", "111"), -- i=1893
      ("0101010001110000", "111"), -- i=1894
      ("0100010001110000", "111"), -- i=1895
      ("1000010001110100", "111"), -- i=1896
      ("1001010001110100", "111"), -- i=1897
      ("1010010001110100", "111"), -- i=1898
      ("1011010001110100", "111"), -- i=1899
      ("0101010001110000", "111"), -- i=1900
      ("0100010001110000", "111"), -- i=1901
      ("1000010001110101", "111"), -- i=1902
      ("1001010001110101", "111"), -- i=1903
      ("1010010001110101", "111"), -- i=1904
      ("1011010001110101", "111"), -- i=1905
      ("0101010001110000", "111"), -- i=1906
      ("0100010001110000", "111"), -- i=1907
      ("1000010001110110", "111"), -- i=1908
      ("1001010001110110", "111"), -- i=1909
      ("1010010001110110", "111"), -- i=1910
      ("1011010001110110", "111"), -- i=1911
      ("0101010001110000", "111"), -- i=1912
      ("0100010001110000", "111"), -- i=1913
      ("1000010001110111", "111"), -- i=1914
      ("1001010001110111", "111"), -- i=1915
      ("1010010001110111", "111"), -- i=1916
      ("1011010001110111", "111"), -- i=1917
      ("0101010001110000", "111"), -- i=1918
      ("0100010001110000", "111"), -- i=1919
      ("1000010100000000", "000"), -- i=1920
      ("1001010100000000", "000"), -- i=1921
      ("1010010100000000", "000"), -- i=1922
      ("1011010100000000", "000"), -- i=1923
      ("0101010100000000", "000"), -- i=1924
      ("0100010100000000", "000"), -- i=1925
      ("1000010100000001", "000"), -- i=1926
      ("1001010100000001", "000"), -- i=1927
      ("1010010100000001", "000"), -- i=1928
      ("1011010100000001", "000"), -- i=1929
      ("0101010100000000", "000"), -- i=1930
      ("0100010100000000", "000"), -- i=1931
      ("1000010100000010", "000"), -- i=1932
      ("1001010100000010", "000"), -- i=1933
      ("1010010100000010", "000"), -- i=1934
      ("1011010100000010", "000"), -- i=1935
      ("0101010100000000", "000"), -- i=1936
      ("0100010100000000", "000"), -- i=1937
      ("1000010100000011", "000"), -- i=1938
      ("1001010100000011", "000"), -- i=1939
      ("1010010100000011", "000"), -- i=1940
      ("1011010100000011", "000"), -- i=1941
      ("0101010100000000", "000"), -- i=1942
      ("0100010100000000", "000"), -- i=1943
      ("1000010100000100", "000"), -- i=1944
      ("1001010100000100", "000"), -- i=1945
      ("1010010100000100", "000"), -- i=1946
      ("1011010100000100", "000"), -- i=1947
      ("0101010100000000", "000"), -- i=1948
      ("0100010100000000", "000"), -- i=1949
      ("1000010100000101", "000"), -- i=1950
      ("1001010100000101", "000"), -- i=1951
      ("1010010100000101", "000"), -- i=1952
      ("1011010100000101", "000"), -- i=1953
      ("0101010100000000", "000"), -- i=1954
      ("0100010100000000", "000"), -- i=1955
      ("1000010100000110", "000"), -- i=1956
      ("1001010100000110", "000"), -- i=1957
      ("1010010100000110", "000"), -- i=1958
      ("1011010100000110", "000"), -- i=1959
      ("0101010100000000", "000"), -- i=1960
      ("0100010100000000", "000"), -- i=1961
      ("1000010100000111", "000"), -- i=1962
      ("1001010100000111", "000"), -- i=1963
      ("1010010100000111", "000"), -- i=1964
      ("1011010100000111", "000"), -- i=1965
      ("0101010100000000", "000"), -- i=1966
      ("0100010100000000", "000"), -- i=1967
      ("1000010100010000", "001"), -- i=1968
      ("1001010100010000", "001"), -- i=1969
      ("1010010100010000", "001"), -- i=1970
      ("1011010100010000", "001"), -- i=1971
      ("0101010100010000", "001"), -- i=1972
      ("0100010100010000", "001"), -- i=1973
      ("1000010100010001", "001"), -- i=1974
      ("1001010100010001", "001"), -- i=1975
      ("1010010100010001", "001"), -- i=1976
      ("1011010100010001", "001"), -- i=1977
      ("0101010100010000", "001"), -- i=1978
      ("0100010100010000", "001"), -- i=1979
      ("1000010100010010", "001"), -- i=1980
      ("1001010100010010", "001"), -- i=1981
      ("1010010100010010", "001"), -- i=1982
      ("1011010100010010", "001"), -- i=1983
      ("0101010100010000", "001"), -- i=1984
      ("0100010100010000", "001"), -- i=1985
      ("1000010100010011", "001"), -- i=1986
      ("1001010100010011", "001"), -- i=1987
      ("1010010100010011", "001"), -- i=1988
      ("1011010100010011", "001"), -- i=1989
      ("0101010100010000", "001"), -- i=1990
      ("0100010100010000", "001"), -- i=1991
      ("1000010100010100", "001"), -- i=1992
      ("1001010100010100", "001"), -- i=1993
      ("1010010100010100", "001"), -- i=1994
      ("1011010100010100", "001"), -- i=1995
      ("0101010100010000", "001"), -- i=1996
      ("0100010100010000", "001"), -- i=1997
      ("1000010100010101", "001"), -- i=1998
      ("1001010100010101", "001"), -- i=1999
      ("1010010100010101", "001"), -- i=2000
      ("1011010100010101", "001"), -- i=2001
      ("0101010100010000", "001"), -- i=2002
      ("0100010100010000", "001"), -- i=2003
      ("1000010100010110", "001"), -- i=2004
      ("1001010100010110", "001"), -- i=2005
      ("1010010100010110", "001"), -- i=2006
      ("1011010100010110", "001"), -- i=2007
      ("0101010100010000", "001"), -- i=2008
      ("0100010100010000", "001"), -- i=2009
      ("1000010100010111", "001"), -- i=2010
      ("1001010100010111", "001"), -- i=2011
      ("1010010100010111", "001"), -- i=2012
      ("1011010100010111", "001"), -- i=2013
      ("0101010100010000", "001"), -- i=2014
      ("0100010100010000", "001"), -- i=2015
      ("1000010100100000", "010"), -- i=2016
      ("1001010100100000", "010"), -- i=2017
      ("1010010100100000", "010"), -- i=2018
      ("1011010100100000", "010"), -- i=2019
      ("0101010100100000", "010"), -- i=2020
      ("0100010100100000", "010"), -- i=2021
      ("1000010100100001", "010"), -- i=2022
      ("1001010100100001", "010"), -- i=2023
      ("1010010100100001", "010"), -- i=2024
      ("1011010100100001", "010"), -- i=2025
      ("0101010100100000", "010"), -- i=2026
      ("0100010100100000", "010"), -- i=2027
      ("1000010100100010", "010"), -- i=2028
      ("1001010100100010", "010"), -- i=2029
      ("1010010100100010", "010"), -- i=2030
      ("1011010100100010", "010"), -- i=2031
      ("0101010100100000", "010"), -- i=2032
      ("0100010100100000", "010"), -- i=2033
      ("1000010100100011", "010"), -- i=2034
      ("1001010100100011", "010"), -- i=2035
      ("1010010100100011", "010"), -- i=2036
      ("1011010100100011", "010"), -- i=2037
      ("0101010100100000", "010"), -- i=2038
      ("0100010100100000", "010"), -- i=2039
      ("1000010100100100", "010"), -- i=2040
      ("1001010100100100", "010"), -- i=2041
      ("1010010100100100", "010"), -- i=2042
      ("1011010100100100", "010"), -- i=2043
      ("0101010100100000", "010"), -- i=2044
      ("0100010100100000", "010"), -- i=2045
      ("1000010100100101", "010"), -- i=2046
      ("1001010100100101", "010"), -- i=2047
      ("1010010100100101", "010"), -- i=2048
      ("1011010100100101", "010"), -- i=2049
      ("0101010100100000", "010"), -- i=2050
      ("0100010100100000", "010"), -- i=2051
      ("1000010100100110", "010"), -- i=2052
      ("1001010100100110", "010"), -- i=2053
      ("1010010100100110", "010"), -- i=2054
      ("1011010100100110", "010"), -- i=2055
      ("0101010100100000", "010"), -- i=2056
      ("0100010100100000", "010"), -- i=2057
      ("1000010100100111", "010"), -- i=2058
      ("1001010100100111", "010"), -- i=2059
      ("1010010100100111", "010"), -- i=2060
      ("1011010100100111", "010"), -- i=2061
      ("0101010100100000", "010"), -- i=2062
      ("0100010100100000", "010"), -- i=2063
      ("1000010100110000", "011"), -- i=2064
      ("1001010100110000", "011"), -- i=2065
      ("1010010100110000", "011"), -- i=2066
      ("1011010100110000", "011"), -- i=2067
      ("0101010100110000", "011"), -- i=2068
      ("0100010100110000", "011"), -- i=2069
      ("1000010100110001", "011"), -- i=2070
      ("1001010100110001", "011"), -- i=2071
      ("1010010100110001", "011"), -- i=2072
      ("1011010100110001", "011"), -- i=2073
      ("0101010100110000", "011"), -- i=2074
      ("0100010100110000", "011"), -- i=2075
      ("1000010100110010", "011"), -- i=2076
      ("1001010100110010", "011"), -- i=2077
      ("1010010100110010", "011"), -- i=2078
      ("1011010100110010", "011"), -- i=2079
      ("0101010100110000", "011"), -- i=2080
      ("0100010100110000", "011"), -- i=2081
      ("1000010100110011", "011"), -- i=2082
      ("1001010100110011", "011"), -- i=2083
      ("1010010100110011", "011"), -- i=2084
      ("1011010100110011", "011"), -- i=2085
      ("0101010100110000", "011"), -- i=2086
      ("0100010100110000", "011"), -- i=2087
      ("1000010100110100", "011"), -- i=2088
      ("1001010100110100", "011"), -- i=2089
      ("1010010100110100", "011"), -- i=2090
      ("1011010100110100", "011"), -- i=2091
      ("0101010100110000", "011"), -- i=2092
      ("0100010100110000", "011"), -- i=2093
      ("1000010100110101", "011"), -- i=2094
      ("1001010100110101", "011"), -- i=2095
      ("1010010100110101", "011"), -- i=2096
      ("1011010100110101", "011"), -- i=2097
      ("0101010100110000", "011"), -- i=2098
      ("0100010100110000", "011"), -- i=2099
      ("1000010100110110", "011"), -- i=2100
      ("1001010100110110", "011"), -- i=2101
      ("1010010100110110", "011"), -- i=2102
      ("1011010100110110", "011"), -- i=2103
      ("0101010100110000", "011"), -- i=2104
      ("0100010100110000", "011"), -- i=2105
      ("1000010100110111", "011"), -- i=2106
      ("1001010100110111", "011"), -- i=2107
      ("1010010100110111", "011"), -- i=2108
      ("1011010100110111", "011"), -- i=2109
      ("0101010100110000", "011"), -- i=2110
      ("0100010100110000", "011"), -- i=2111
      ("1000010101000000", "100"), -- i=2112
      ("1001010101000000", "100"), -- i=2113
      ("1010010101000000", "100"), -- i=2114
      ("1011010101000000", "100"), -- i=2115
      ("0101010101000000", "100"), -- i=2116
      ("0100010101000000", "100"), -- i=2117
      ("1000010101000001", "100"), -- i=2118
      ("1001010101000001", "100"), -- i=2119
      ("1010010101000001", "100"), -- i=2120
      ("1011010101000001", "100"), -- i=2121
      ("0101010101000000", "100"), -- i=2122
      ("0100010101000000", "100"), -- i=2123
      ("1000010101000010", "100"), -- i=2124
      ("1001010101000010", "100"), -- i=2125
      ("1010010101000010", "100"), -- i=2126
      ("1011010101000010", "100"), -- i=2127
      ("0101010101000000", "100"), -- i=2128
      ("0100010101000000", "100"), -- i=2129
      ("1000010101000011", "100"), -- i=2130
      ("1001010101000011", "100"), -- i=2131
      ("1010010101000011", "100"), -- i=2132
      ("1011010101000011", "100"), -- i=2133
      ("0101010101000000", "100"), -- i=2134
      ("0100010101000000", "100"), -- i=2135
      ("1000010101000100", "100"), -- i=2136
      ("1001010101000100", "100"), -- i=2137
      ("1010010101000100", "100"), -- i=2138
      ("1011010101000100", "100"), -- i=2139
      ("0101010101000000", "100"), -- i=2140
      ("0100010101000000", "100"), -- i=2141
      ("1000010101000101", "100"), -- i=2142
      ("1001010101000101", "100"), -- i=2143
      ("1010010101000101", "100"), -- i=2144
      ("1011010101000101", "100"), -- i=2145
      ("0101010101000000", "100"), -- i=2146
      ("0100010101000000", "100"), -- i=2147
      ("1000010101000110", "100"), -- i=2148
      ("1001010101000110", "100"), -- i=2149
      ("1010010101000110", "100"), -- i=2150
      ("1011010101000110", "100"), -- i=2151
      ("0101010101000000", "100"), -- i=2152
      ("0100010101000000", "100"), -- i=2153
      ("1000010101000111", "100"), -- i=2154
      ("1001010101000111", "100"), -- i=2155
      ("1010010101000111", "100"), -- i=2156
      ("1011010101000111", "100"), -- i=2157
      ("0101010101000000", "100"), -- i=2158
      ("0100010101000000", "100"), -- i=2159
      ("1000010101010000", "101"), -- i=2160
      ("1001010101010000", "101"), -- i=2161
      ("1010010101010000", "101"), -- i=2162
      ("1011010101010000", "101"), -- i=2163
      ("0101010101010000", "101"), -- i=2164
      ("0100010101010000", "101"), -- i=2165
      ("1000010101010001", "101"), -- i=2166
      ("1001010101010001", "101"), -- i=2167
      ("1010010101010001", "101"), -- i=2168
      ("1011010101010001", "101"), -- i=2169
      ("0101010101010000", "101"), -- i=2170
      ("0100010101010000", "101"), -- i=2171
      ("1000010101010010", "101"), -- i=2172
      ("1001010101010010", "101"), -- i=2173
      ("1010010101010010", "101"), -- i=2174
      ("1011010101010010", "101"), -- i=2175
      ("0101010101010000", "101"), -- i=2176
      ("0100010101010000", "101"), -- i=2177
      ("1000010101010011", "101"), -- i=2178
      ("1001010101010011", "101"), -- i=2179
      ("1010010101010011", "101"), -- i=2180
      ("1011010101010011", "101"), -- i=2181
      ("0101010101010000", "101"), -- i=2182
      ("0100010101010000", "101"), -- i=2183
      ("1000010101010100", "101"), -- i=2184
      ("1001010101010100", "101"), -- i=2185
      ("1010010101010100", "101"), -- i=2186
      ("1011010101010100", "101"), -- i=2187
      ("0101010101010000", "101"), -- i=2188
      ("0100010101010000", "101"), -- i=2189
      ("1000010101010101", "101"), -- i=2190
      ("1001010101010101", "101"), -- i=2191
      ("1010010101010101", "101"), -- i=2192
      ("1011010101010101", "101"), -- i=2193
      ("0101010101010000", "101"), -- i=2194
      ("0100010101010000", "101"), -- i=2195
      ("1000010101010110", "101"), -- i=2196
      ("1001010101010110", "101"), -- i=2197
      ("1010010101010110", "101"), -- i=2198
      ("1011010101010110", "101"), -- i=2199
      ("0101010101010000", "101"), -- i=2200
      ("0100010101010000", "101"), -- i=2201
      ("1000010101010111", "101"), -- i=2202
      ("1001010101010111", "101"), -- i=2203
      ("1010010101010111", "101"), -- i=2204
      ("1011010101010111", "101"), -- i=2205
      ("0101010101010000", "101"), -- i=2206
      ("0100010101010000", "101"), -- i=2207
      ("1000010101100000", "110"), -- i=2208
      ("1001010101100000", "110"), -- i=2209
      ("1010010101100000", "110"), -- i=2210
      ("1011010101100000", "110"), -- i=2211
      ("0101010101100000", "110"), -- i=2212
      ("0100010101100000", "110"), -- i=2213
      ("1000010101100001", "110"), -- i=2214
      ("1001010101100001", "110"), -- i=2215
      ("1010010101100001", "110"), -- i=2216
      ("1011010101100001", "110"), -- i=2217
      ("0101010101100000", "110"), -- i=2218
      ("0100010101100000", "110"), -- i=2219
      ("1000010101100010", "110"), -- i=2220
      ("1001010101100010", "110"), -- i=2221
      ("1010010101100010", "110"), -- i=2222
      ("1011010101100010", "110"), -- i=2223
      ("0101010101100000", "110"), -- i=2224
      ("0100010101100000", "110"), -- i=2225
      ("1000010101100011", "110"), -- i=2226
      ("1001010101100011", "110"), -- i=2227
      ("1010010101100011", "110"), -- i=2228
      ("1011010101100011", "110"), -- i=2229
      ("0101010101100000", "110"), -- i=2230
      ("0100010101100000", "110"), -- i=2231
      ("1000010101100100", "110"), -- i=2232
      ("1001010101100100", "110"), -- i=2233
      ("1010010101100100", "110"), -- i=2234
      ("1011010101100100", "110"), -- i=2235
      ("0101010101100000", "110"), -- i=2236
      ("0100010101100000", "110"), -- i=2237
      ("1000010101100101", "110"), -- i=2238
      ("1001010101100101", "110"), -- i=2239
      ("1010010101100101", "110"), -- i=2240
      ("1011010101100101", "110"), -- i=2241
      ("0101010101100000", "110"), -- i=2242
      ("0100010101100000", "110"), -- i=2243
      ("1000010101100110", "110"), -- i=2244
      ("1001010101100110", "110"), -- i=2245
      ("1010010101100110", "110"), -- i=2246
      ("1011010101100110", "110"), -- i=2247
      ("0101010101100000", "110"), -- i=2248
      ("0100010101100000", "110"), -- i=2249
      ("1000010101100111", "110"), -- i=2250
      ("1001010101100111", "110"), -- i=2251
      ("1010010101100111", "110"), -- i=2252
      ("1011010101100111", "110"), -- i=2253
      ("0101010101100000", "110"), -- i=2254
      ("0100010101100000", "110"), -- i=2255
      ("1000010101110000", "111"), -- i=2256
      ("1001010101110000", "111"), -- i=2257
      ("1010010101110000", "111"), -- i=2258
      ("1011010101110000", "111"), -- i=2259
      ("0101010101110000", "111"), -- i=2260
      ("0100010101110000", "111"), -- i=2261
      ("1000010101110001", "111"), -- i=2262
      ("1001010101110001", "111"), -- i=2263
      ("1010010101110001", "111"), -- i=2264
      ("1011010101110001", "111"), -- i=2265
      ("0101010101110000", "111"), -- i=2266
      ("0100010101110000", "111"), -- i=2267
      ("1000010101110010", "111"), -- i=2268
      ("1001010101110010", "111"), -- i=2269
      ("1010010101110010", "111"), -- i=2270
      ("1011010101110010", "111"), -- i=2271
      ("0101010101110000", "111"), -- i=2272
      ("0100010101110000", "111"), -- i=2273
      ("1000010101110011", "111"), -- i=2274
      ("1001010101110011", "111"), -- i=2275
      ("1010010101110011", "111"), -- i=2276
      ("1011010101110011", "111"), -- i=2277
      ("0101010101110000", "111"), -- i=2278
      ("0100010101110000", "111"), -- i=2279
      ("1000010101110100", "111"), -- i=2280
      ("1001010101110100", "111"), -- i=2281
      ("1010010101110100", "111"), -- i=2282
      ("1011010101110100", "111"), -- i=2283
      ("0101010101110000", "111"), -- i=2284
      ("0100010101110000", "111"), -- i=2285
      ("1000010101110101", "111"), -- i=2286
      ("1001010101110101", "111"), -- i=2287
      ("1010010101110101", "111"), -- i=2288
      ("1011010101110101", "111"), -- i=2289
      ("0101010101110000", "111"), -- i=2290
      ("0100010101110000", "111"), -- i=2291
      ("1000010101110110", "111"), -- i=2292
      ("1001010101110110", "111"), -- i=2293
      ("1010010101110110", "111"), -- i=2294
      ("1011010101110110", "111"), -- i=2295
      ("0101010101110000", "111"), -- i=2296
      ("0100010101110000", "111"), -- i=2297
      ("1000010101110111", "111"), -- i=2298
      ("1001010101110111", "111"), -- i=2299
      ("1010010101110111", "111"), -- i=2300
      ("1011010101110111", "111"), -- i=2301
      ("0101010101110000", "111"), -- i=2302
      ("0100010101110000", "111"), -- i=2303
      ("1000011000000000", "000"), -- i=2304
      ("1001011000000000", "000"), -- i=2305
      ("1010011000000000", "000"), -- i=2306
      ("1011011000000000", "000"), -- i=2307
      ("0101011000000000", "000"), -- i=2308
      ("0100011000000000", "000"), -- i=2309
      ("1000011000000001", "000"), -- i=2310
      ("1001011000000001", "000"), -- i=2311
      ("1010011000000001", "000"), -- i=2312
      ("1011011000000001", "000"), -- i=2313
      ("0101011000000000", "000"), -- i=2314
      ("0100011000000000", "000"), -- i=2315
      ("1000011000000010", "000"), -- i=2316
      ("1001011000000010", "000"), -- i=2317
      ("1010011000000010", "000"), -- i=2318
      ("1011011000000010", "000"), -- i=2319
      ("0101011000000000", "000"), -- i=2320
      ("0100011000000000", "000"), -- i=2321
      ("1000011000000011", "000"), -- i=2322
      ("1001011000000011", "000"), -- i=2323
      ("1010011000000011", "000"), -- i=2324
      ("1011011000000011", "000"), -- i=2325
      ("0101011000000000", "000"), -- i=2326
      ("0100011000000000", "000"), -- i=2327
      ("1000011000000100", "000"), -- i=2328
      ("1001011000000100", "000"), -- i=2329
      ("1010011000000100", "000"), -- i=2330
      ("1011011000000100", "000"), -- i=2331
      ("0101011000000000", "000"), -- i=2332
      ("0100011000000000", "000"), -- i=2333
      ("1000011000000101", "000"), -- i=2334
      ("1001011000000101", "000"), -- i=2335
      ("1010011000000101", "000"), -- i=2336
      ("1011011000000101", "000"), -- i=2337
      ("0101011000000000", "000"), -- i=2338
      ("0100011000000000", "000"), -- i=2339
      ("1000011000000110", "000"), -- i=2340
      ("1001011000000110", "000"), -- i=2341
      ("1010011000000110", "000"), -- i=2342
      ("1011011000000110", "000"), -- i=2343
      ("0101011000000000", "000"), -- i=2344
      ("0100011000000000", "000"), -- i=2345
      ("1000011000000111", "000"), -- i=2346
      ("1001011000000111", "000"), -- i=2347
      ("1010011000000111", "000"), -- i=2348
      ("1011011000000111", "000"), -- i=2349
      ("0101011000000000", "000"), -- i=2350
      ("0100011000000000", "000"), -- i=2351
      ("1000011000010000", "001"), -- i=2352
      ("1001011000010000", "001"), -- i=2353
      ("1010011000010000", "001"), -- i=2354
      ("1011011000010000", "001"), -- i=2355
      ("0101011000010000", "001"), -- i=2356
      ("0100011000010000", "001"), -- i=2357
      ("1000011000010001", "001"), -- i=2358
      ("1001011000010001", "001"), -- i=2359
      ("1010011000010001", "001"), -- i=2360
      ("1011011000010001", "001"), -- i=2361
      ("0101011000010000", "001"), -- i=2362
      ("0100011000010000", "001"), -- i=2363
      ("1000011000010010", "001"), -- i=2364
      ("1001011000010010", "001"), -- i=2365
      ("1010011000010010", "001"), -- i=2366
      ("1011011000010010", "001"), -- i=2367
      ("0101011000010000", "001"), -- i=2368
      ("0100011000010000", "001"), -- i=2369
      ("1000011000010011", "001"), -- i=2370
      ("1001011000010011", "001"), -- i=2371
      ("1010011000010011", "001"), -- i=2372
      ("1011011000010011", "001"), -- i=2373
      ("0101011000010000", "001"), -- i=2374
      ("0100011000010000", "001"), -- i=2375
      ("1000011000010100", "001"), -- i=2376
      ("1001011000010100", "001"), -- i=2377
      ("1010011000010100", "001"), -- i=2378
      ("1011011000010100", "001"), -- i=2379
      ("0101011000010000", "001"), -- i=2380
      ("0100011000010000", "001"), -- i=2381
      ("1000011000010101", "001"), -- i=2382
      ("1001011000010101", "001"), -- i=2383
      ("1010011000010101", "001"), -- i=2384
      ("1011011000010101", "001"), -- i=2385
      ("0101011000010000", "001"), -- i=2386
      ("0100011000010000", "001"), -- i=2387
      ("1000011000010110", "001"), -- i=2388
      ("1001011000010110", "001"), -- i=2389
      ("1010011000010110", "001"), -- i=2390
      ("1011011000010110", "001"), -- i=2391
      ("0101011000010000", "001"), -- i=2392
      ("0100011000010000", "001"), -- i=2393
      ("1000011000010111", "001"), -- i=2394
      ("1001011000010111", "001"), -- i=2395
      ("1010011000010111", "001"), -- i=2396
      ("1011011000010111", "001"), -- i=2397
      ("0101011000010000", "001"), -- i=2398
      ("0100011000010000", "001"), -- i=2399
      ("1000011000100000", "010"), -- i=2400
      ("1001011000100000", "010"), -- i=2401
      ("1010011000100000", "010"), -- i=2402
      ("1011011000100000", "010"), -- i=2403
      ("0101011000100000", "010"), -- i=2404
      ("0100011000100000", "010"), -- i=2405
      ("1000011000100001", "010"), -- i=2406
      ("1001011000100001", "010"), -- i=2407
      ("1010011000100001", "010"), -- i=2408
      ("1011011000100001", "010"), -- i=2409
      ("0101011000100000", "010"), -- i=2410
      ("0100011000100000", "010"), -- i=2411
      ("1000011000100010", "010"), -- i=2412
      ("1001011000100010", "010"), -- i=2413
      ("1010011000100010", "010"), -- i=2414
      ("1011011000100010", "010"), -- i=2415
      ("0101011000100000", "010"), -- i=2416
      ("0100011000100000", "010"), -- i=2417
      ("1000011000100011", "010"), -- i=2418
      ("1001011000100011", "010"), -- i=2419
      ("1010011000100011", "010"), -- i=2420
      ("1011011000100011", "010"), -- i=2421
      ("0101011000100000", "010"), -- i=2422
      ("0100011000100000", "010"), -- i=2423
      ("1000011000100100", "010"), -- i=2424
      ("1001011000100100", "010"), -- i=2425
      ("1010011000100100", "010"), -- i=2426
      ("1011011000100100", "010"), -- i=2427
      ("0101011000100000", "010"), -- i=2428
      ("0100011000100000", "010"), -- i=2429
      ("1000011000100101", "010"), -- i=2430
      ("1001011000100101", "010"), -- i=2431
      ("1010011000100101", "010"), -- i=2432
      ("1011011000100101", "010"), -- i=2433
      ("0101011000100000", "010"), -- i=2434
      ("0100011000100000", "010"), -- i=2435
      ("1000011000100110", "010"), -- i=2436
      ("1001011000100110", "010"), -- i=2437
      ("1010011000100110", "010"), -- i=2438
      ("1011011000100110", "010"), -- i=2439
      ("0101011000100000", "010"), -- i=2440
      ("0100011000100000", "010"), -- i=2441
      ("1000011000100111", "010"), -- i=2442
      ("1001011000100111", "010"), -- i=2443
      ("1010011000100111", "010"), -- i=2444
      ("1011011000100111", "010"), -- i=2445
      ("0101011000100000", "010"), -- i=2446
      ("0100011000100000", "010"), -- i=2447
      ("1000011000110000", "011"), -- i=2448
      ("1001011000110000", "011"), -- i=2449
      ("1010011000110000", "011"), -- i=2450
      ("1011011000110000", "011"), -- i=2451
      ("0101011000110000", "011"), -- i=2452
      ("0100011000110000", "011"), -- i=2453
      ("1000011000110001", "011"), -- i=2454
      ("1001011000110001", "011"), -- i=2455
      ("1010011000110001", "011"), -- i=2456
      ("1011011000110001", "011"), -- i=2457
      ("0101011000110000", "011"), -- i=2458
      ("0100011000110000", "011"), -- i=2459
      ("1000011000110010", "011"), -- i=2460
      ("1001011000110010", "011"), -- i=2461
      ("1010011000110010", "011"), -- i=2462
      ("1011011000110010", "011"), -- i=2463
      ("0101011000110000", "011"), -- i=2464
      ("0100011000110000", "011"), -- i=2465
      ("1000011000110011", "011"), -- i=2466
      ("1001011000110011", "011"), -- i=2467
      ("1010011000110011", "011"), -- i=2468
      ("1011011000110011", "011"), -- i=2469
      ("0101011000110000", "011"), -- i=2470
      ("0100011000110000", "011"), -- i=2471
      ("1000011000110100", "011"), -- i=2472
      ("1001011000110100", "011"), -- i=2473
      ("1010011000110100", "011"), -- i=2474
      ("1011011000110100", "011"), -- i=2475
      ("0101011000110000", "011"), -- i=2476
      ("0100011000110000", "011"), -- i=2477
      ("1000011000110101", "011"), -- i=2478
      ("1001011000110101", "011"), -- i=2479
      ("1010011000110101", "011"), -- i=2480
      ("1011011000110101", "011"), -- i=2481
      ("0101011000110000", "011"), -- i=2482
      ("0100011000110000", "011"), -- i=2483
      ("1000011000110110", "011"), -- i=2484
      ("1001011000110110", "011"), -- i=2485
      ("1010011000110110", "011"), -- i=2486
      ("1011011000110110", "011"), -- i=2487
      ("0101011000110000", "011"), -- i=2488
      ("0100011000110000", "011"), -- i=2489
      ("1000011000110111", "011"), -- i=2490
      ("1001011000110111", "011"), -- i=2491
      ("1010011000110111", "011"), -- i=2492
      ("1011011000110111", "011"), -- i=2493
      ("0101011000110000", "011"), -- i=2494
      ("0100011000110000", "011"), -- i=2495
      ("1000011001000000", "100"), -- i=2496
      ("1001011001000000", "100"), -- i=2497
      ("1010011001000000", "100"), -- i=2498
      ("1011011001000000", "100"), -- i=2499
      ("0101011001000000", "100"), -- i=2500
      ("0100011001000000", "100"), -- i=2501
      ("1000011001000001", "100"), -- i=2502
      ("1001011001000001", "100"), -- i=2503
      ("1010011001000001", "100"), -- i=2504
      ("1011011001000001", "100"), -- i=2505
      ("0101011001000000", "100"), -- i=2506
      ("0100011001000000", "100"), -- i=2507
      ("1000011001000010", "100"), -- i=2508
      ("1001011001000010", "100"), -- i=2509
      ("1010011001000010", "100"), -- i=2510
      ("1011011001000010", "100"), -- i=2511
      ("0101011001000000", "100"), -- i=2512
      ("0100011001000000", "100"), -- i=2513
      ("1000011001000011", "100"), -- i=2514
      ("1001011001000011", "100"), -- i=2515
      ("1010011001000011", "100"), -- i=2516
      ("1011011001000011", "100"), -- i=2517
      ("0101011001000000", "100"), -- i=2518
      ("0100011001000000", "100"), -- i=2519
      ("1000011001000100", "100"), -- i=2520
      ("1001011001000100", "100"), -- i=2521
      ("1010011001000100", "100"), -- i=2522
      ("1011011001000100", "100"), -- i=2523
      ("0101011001000000", "100"), -- i=2524
      ("0100011001000000", "100"), -- i=2525
      ("1000011001000101", "100"), -- i=2526
      ("1001011001000101", "100"), -- i=2527
      ("1010011001000101", "100"), -- i=2528
      ("1011011001000101", "100"), -- i=2529
      ("0101011001000000", "100"), -- i=2530
      ("0100011001000000", "100"), -- i=2531
      ("1000011001000110", "100"), -- i=2532
      ("1001011001000110", "100"), -- i=2533
      ("1010011001000110", "100"), -- i=2534
      ("1011011001000110", "100"), -- i=2535
      ("0101011001000000", "100"), -- i=2536
      ("0100011001000000", "100"), -- i=2537
      ("1000011001000111", "100"), -- i=2538
      ("1001011001000111", "100"), -- i=2539
      ("1010011001000111", "100"), -- i=2540
      ("1011011001000111", "100"), -- i=2541
      ("0101011001000000", "100"), -- i=2542
      ("0100011001000000", "100"), -- i=2543
      ("1000011001010000", "101"), -- i=2544
      ("1001011001010000", "101"), -- i=2545
      ("1010011001010000", "101"), -- i=2546
      ("1011011001010000", "101"), -- i=2547
      ("0101011001010000", "101"), -- i=2548
      ("0100011001010000", "101"), -- i=2549
      ("1000011001010001", "101"), -- i=2550
      ("1001011001010001", "101"), -- i=2551
      ("1010011001010001", "101"), -- i=2552
      ("1011011001010001", "101"), -- i=2553
      ("0101011001010000", "101"), -- i=2554
      ("0100011001010000", "101"), -- i=2555
      ("1000011001010010", "101"), -- i=2556
      ("1001011001010010", "101"), -- i=2557
      ("1010011001010010", "101"), -- i=2558
      ("1011011001010010", "101"), -- i=2559
      ("0101011001010000", "101"), -- i=2560
      ("0100011001010000", "101"), -- i=2561
      ("1000011001010011", "101"), -- i=2562
      ("1001011001010011", "101"), -- i=2563
      ("1010011001010011", "101"), -- i=2564
      ("1011011001010011", "101"), -- i=2565
      ("0101011001010000", "101"), -- i=2566
      ("0100011001010000", "101"), -- i=2567
      ("1000011001010100", "101"), -- i=2568
      ("1001011001010100", "101"), -- i=2569
      ("1010011001010100", "101"), -- i=2570
      ("1011011001010100", "101"), -- i=2571
      ("0101011001010000", "101"), -- i=2572
      ("0100011001010000", "101"), -- i=2573
      ("1000011001010101", "101"), -- i=2574
      ("1001011001010101", "101"), -- i=2575
      ("1010011001010101", "101"), -- i=2576
      ("1011011001010101", "101"), -- i=2577
      ("0101011001010000", "101"), -- i=2578
      ("0100011001010000", "101"), -- i=2579
      ("1000011001010110", "101"), -- i=2580
      ("1001011001010110", "101"), -- i=2581
      ("1010011001010110", "101"), -- i=2582
      ("1011011001010110", "101"), -- i=2583
      ("0101011001010000", "101"), -- i=2584
      ("0100011001010000", "101"), -- i=2585
      ("1000011001010111", "101"), -- i=2586
      ("1001011001010111", "101"), -- i=2587
      ("1010011001010111", "101"), -- i=2588
      ("1011011001010111", "101"), -- i=2589
      ("0101011001010000", "101"), -- i=2590
      ("0100011001010000", "101"), -- i=2591
      ("1000011001100000", "110"), -- i=2592
      ("1001011001100000", "110"), -- i=2593
      ("1010011001100000", "110"), -- i=2594
      ("1011011001100000", "110"), -- i=2595
      ("0101011001100000", "110"), -- i=2596
      ("0100011001100000", "110"), -- i=2597
      ("1000011001100001", "110"), -- i=2598
      ("1001011001100001", "110"), -- i=2599
      ("1010011001100001", "110"), -- i=2600
      ("1011011001100001", "110"), -- i=2601
      ("0101011001100000", "110"), -- i=2602
      ("0100011001100000", "110"), -- i=2603
      ("1000011001100010", "110"), -- i=2604
      ("1001011001100010", "110"), -- i=2605
      ("1010011001100010", "110"), -- i=2606
      ("1011011001100010", "110"), -- i=2607
      ("0101011001100000", "110"), -- i=2608
      ("0100011001100000", "110"), -- i=2609
      ("1000011001100011", "110"), -- i=2610
      ("1001011001100011", "110"), -- i=2611
      ("1010011001100011", "110"), -- i=2612
      ("1011011001100011", "110"), -- i=2613
      ("0101011001100000", "110"), -- i=2614
      ("0100011001100000", "110"), -- i=2615
      ("1000011001100100", "110"), -- i=2616
      ("1001011001100100", "110"), -- i=2617
      ("1010011001100100", "110"), -- i=2618
      ("1011011001100100", "110"), -- i=2619
      ("0101011001100000", "110"), -- i=2620
      ("0100011001100000", "110"), -- i=2621
      ("1000011001100101", "110"), -- i=2622
      ("1001011001100101", "110"), -- i=2623
      ("1010011001100101", "110"), -- i=2624
      ("1011011001100101", "110"), -- i=2625
      ("0101011001100000", "110"), -- i=2626
      ("0100011001100000", "110"), -- i=2627
      ("1000011001100110", "110"), -- i=2628
      ("1001011001100110", "110"), -- i=2629
      ("1010011001100110", "110"), -- i=2630
      ("1011011001100110", "110"), -- i=2631
      ("0101011001100000", "110"), -- i=2632
      ("0100011001100000", "110"), -- i=2633
      ("1000011001100111", "110"), -- i=2634
      ("1001011001100111", "110"), -- i=2635
      ("1010011001100111", "110"), -- i=2636
      ("1011011001100111", "110"), -- i=2637
      ("0101011001100000", "110"), -- i=2638
      ("0100011001100000", "110"), -- i=2639
      ("1000011001110000", "111"), -- i=2640
      ("1001011001110000", "111"), -- i=2641
      ("1010011001110000", "111"), -- i=2642
      ("1011011001110000", "111"), -- i=2643
      ("0101011001110000", "111"), -- i=2644
      ("0100011001110000", "111"), -- i=2645
      ("1000011001110001", "111"), -- i=2646
      ("1001011001110001", "111"), -- i=2647
      ("1010011001110001", "111"), -- i=2648
      ("1011011001110001", "111"), -- i=2649
      ("0101011001110000", "111"), -- i=2650
      ("0100011001110000", "111"), -- i=2651
      ("1000011001110010", "111"), -- i=2652
      ("1001011001110010", "111"), -- i=2653
      ("1010011001110010", "111"), -- i=2654
      ("1011011001110010", "111"), -- i=2655
      ("0101011001110000", "111"), -- i=2656
      ("0100011001110000", "111"), -- i=2657
      ("1000011001110011", "111"), -- i=2658
      ("1001011001110011", "111"), -- i=2659
      ("1010011001110011", "111"), -- i=2660
      ("1011011001110011", "111"), -- i=2661
      ("0101011001110000", "111"), -- i=2662
      ("0100011001110000", "111"), -- i=2663
      ("1000011001110100", "111"), -- i=2664
      ("1001011001110100", "111"), -- i=2665
      ("1010011001110100", "111"), -- i=2666
      ("1011011001110100", "111"), -- i=2667
      ("0101011001110000", "111"), -- i=2668
      ("0100011001110000", "111"), -- i=2669
      ("1000011001110101", "111"), -- i=2670
      ("1001011001110101", "111"), -- i=2671
      ("1010011001110101", "111"), -- i=2672
      ("1011011001110101", "111"), -- i=2673
      ("0101011001110000", "111"), -- i=2674
      ("0100011001110000", "111"), -- i=2675
      ("1000011001110110", "111"), -- i=2676
      ("1001011001110110", "111"), -- i=2677
      ("1010011001110110", "111"), -- i=2678
      ("1011011001110110", "111"), -- i=2679
      ("0101011001110000", "111"), -- i=2680
      ("0100011001110000", "111"), -- i=2681
      ("1000011001110111", "111"), -- i=2682
      ("1001011001110111", "111"), -- i=2683
      ("1010011001110111", "111"), -- i=2684
      ("1011011001110111", "111"), -- i=2685
      ("0101011001110000", "111"), -- i=2686
      ("0100011001110000", "111"), -- i=2687
      ("1000011100000000", "000"), -- i=2688
      ("1001011100000000", "000"), -- i=2689
      ("1010011100000000", "000"), -- i=2690
      ("1011011100000000", "000"), -- i=2691
      ("0101011100000000", "000"), -- i=2692
      ("0100011100000000", "000"), -- i=2693
      ("1000011100000001", "000"), -- i=2694
      ("1001011100000001", "000"), -- i=2695
      ("1010011100000001", "000"), -- i=2696
      ("1011011100000001", "000"), -- i=2697
      ("0101011100000000", "000"), -- i=2698
      ("0100011100000000", "000"), -- i=2699
      ("1000011100000010", "000"), -- i=2700
      ("1001011100000010", "000"), -- i=2701
      ("1010011100000010", "000"), -- i=2702
      ("1011011100000010", "000"), -- i=2703
      ("0101011100000000", "000"), -- i=2704
      ("0100011100000000", "000"), -- i=2705
      ("1000011100000011", "000"), -- i=2706
      ("1001011100000011", "000"), -- i=2707
      ("1010011100000011", "000"), -- i=2708
      ("1011011100000011", "000"), -- i=2709
      ("0101011100000000", "000"), -- i=2710
      ("0100011100000000", "000"), -- i=2711
      ("1000011100000100", "000"), -- i=2712
      ("1001011100000100", "000"), -- i=2713
      ("1010011100000100", "000"), -- i=2714
      ("1011011100000100", "000"), -- i=2715
      ("0101011100000000", "000"), -- i=2716
      ("0100011100000000", "000"), -- i=2717
      ("1000011100000101", "000"), -- i=2718
      ("1001011100000101", "000"), -- i=2719
      ("1010011100000101", "000"), -- i=2720
      ("1011011100000101", "000"), -- i=2721
      ("0101011100000000", "000"), -- i=2722
      ("0100011100000000", "000"), -- i=2723
      ("1000011100000110", "000"), -- i=2724
      ("1001011100000110", "000"), -- i=2725
      ("1010011100000110", "000"), -- i=2726
      ("1011011100000110", "000"), -- i=2727
      ("0101011100000000", "000"), -- i=2728
      ("0100011100000000", "000"), -- i=2729
      ("1000011100000111", "000"), -- i=2730
      ("1001011100000111", "000"), -- i=2731
      ("1010011100000111", "000"), -- i=2732
      ("1011011100000111", "000"), -- i=2733
      ("0101011100000000", "000"), -- i=2734
      ("0100011100000000", "000"), -- i=2735
      ("1000011100010000", "001"), -- i=2736
      ("1001011100010000", "001"), -- i=2737
      ("1010011100010000", "001"), -- i=2738
      ("1011011100010000", "001"), -- i=2739
      ("0101011100010000", "001"), -- i=2740
      ("0100011100010000", "001"), -- i=2741
      ("1000011100010001", "001"), -- i=2742
      ("1001011100010001", "001"), -- i=2743
      ("1010011100010001", "001"), -- i=2744
      ("1011011100010001", "001"), -- i=2745
      ("0101011100010000", "001"), -- i=2746
      ("0100011100010000", "001"), -- i=2747
      ("1000011100010010", "001"), -- i=2748
      ("1001011100010010", "001"), -- i=2749
      ("1010011100010010", "001"), -- i=2750
      ("1011011100010010", "001"), -- i=2751
      ("0101011100010000", "001"), -- i=2752
      ("0100011100010000", "001"), -- i=2753
      ("1000011100010011", "001"), -- i=2754
      ("1001011100010011", "001"), -- i=2755
      ("1010011100010011", "001"), -- i=2756
      ("1011011100010011", "001"), -- i=2757
      ("0101011100010000", "001"), -- i=2758
      ("0100011100010000", "001"), -- i=2759
      ("1000011100010100", "001"), -- i=2760
      ("1001011100010100", "001"), -- i=2761
      ("1010011100010100", "001"), -- i=2762
      ("1011011100010100", "001"), -- i=2763
      ("0101011100010000", "001"), -- i=2764
      ("0100011100010000", "001"), -- i=2765
      ("1000011100010101", "001"), -- i=2766
      ("1001011100010101", "001"), -- i=2767
      ("1010011100010101", "001"), -- i=2768
      ("1011011100010101", "001"), -- i=2769
      ("0101011100010000", "001"), -- i=2770
      ("0100011100010000", "001"), -- i=2771
      ("1000011100010110", "001"), -- i=2772
      ("1001011100010110", "001"), -- i=2773
      ("1010011100010110", "001"), -- i=2774
      ("1011011100010110", "001"), -- i=2775
      ("0101011100010000", "001"), -- i=2776
      ("0100011100010000", "001"), -- i=2777
      ("1000011100010111", "001"), -- i=2778
      ("1001011100010111", "001"), -- i=2779
      ("1010011100010111", "001"), -- i=2780
      ("1011011100010111", "001"), -- i=2781
      ("0101011100010000", "001"), -- i=2782
      ("0100011100010000", "001"), -- i=2783
      ("1000011100100000", "010"), -- i=2784
      ("1001011100100000", "010"), -- i=2785
      ("1010011100100000", "010"), -- i=2786
      ("1011011100100000", "010"), -- i=2787
      ("0101011100100000", "010"), -- i=2788
      ("0100011100100000", "010"), -- i=2789
      ("1000011100100001", "010"), -- i=2790
      ("1001011100100001", "010"), -- i=2791
      ("1010011100100001", "010"), -- i=2792
      ("1011011100100001", "010"), -- i=2793
      ("0101011100100000", "010"), -- i=2794
      ("0100011100100000", "010"), -- i=2795
      ("1000011100100010", "010"), -- i=2796
      ("1001011100100010", "010"), -- i=2797
      ("1010011100100010", "010"), -- i=2798
      ("1011011100100010", "010"), -- i=2799
      ("0101011100100000", "010"), -- i=2800
      ("0100011100100000", "010"), -- i=2801
      ("1000011100100011", "010"), -- i=2802
      ("1001011100100011", "010"), -- i=2803
      ("1010011100100011", "010"), -- i=2804
      ("1011011100100011", "010"), -- i=2805
      ("0101011100100000", "010"), -- i=2806
      ("0100011100100000", "010"), -- i=2807
      ("1000011100100100", "010"), -- i=2808
      ("1001011100100100", "010"), -- i=2809
      ("1010011100100100", "010"), -- i=2810
      ("1011011100100100", "010"), -- i=2811
      ("0101011100100000", "010"), -- i=2812
      ("0100011100100000", "010"), -- i=2813
      ("1000011100100101", "010"), -- i=2814
      ("1001011100100101", "010"), -- i=2815
      ("1010011100100101", "010"), -- i=2816
      ("1011011100100101", "010"), -- i=2817
      ("0101011100100000", "010"), -- i=2818
      ("0100011100100000", "010"), -- i=2819
      ("1000011100100110", "010"), -- i=2820
      ("1001011100100110", "010"), -- i=2821
      ("1010011100100110", "010"), -- i=2822
      ("1011011100100110", "010"), -- i=2823
      ("0101011100100000", "010"), -- i=2824
      ("0100011100100000", "010"), -- i=2825
      ("1000011100100111", "010"), -- i=2826
      ("1001011100100111", "010"), -- i=2827
      ("1010011100100111", "010"), -- i=2828
      ("1011011100100111", "010"), -- i=2829
      ("0101011100100000", "010"), -- i=2830
      ("0100011100100000", "010"), -- i=2831
      ("1000011100110000", "011"), -- i=2832
      ("1001011100110000", "011"), -- i=2833
      ("1010011100110000", "011"), -- i=2834
      ("1011011100110000", "011"), -- i=2835
      ("0101011100110000", "011"), -- i=2836
      ("0100011100110000", "011"), -- i=2837
      ("1000011100110001", "011"), -- i=2838
      ("1001011100110001", "011"), -- i=2839
      ("1010011100110001", "011"), -- i=2840
      ("1011011100110001", "011"), -- i=2841
      ("0101011100110000", "011"), -- i=2842
      ("0100011100110000", "011"), -- i=2843
      ("1000011100110010", "011"), -- i=2844
      ("1001011100110010", "011"), -- i=2845
      ("1010011100110010", "011"), -- i=2846
      ("1011011100110010", "011"), -- i=2847
      ("0101011100110000", "011"), -- i=2848
      ("0100011100110000", "011"), -- i=2849
      ("1000011100110011", "011"), -- i=2850
      ("1001011100110011", "011"), -- i=2851
      ("1010011100110011", "011"), -- i=2852
      ("1011011100110011", "011"), -- i=2853
      ("0101011100110000", "011"), -- i=2854
      ("0100011100110000", "011"), -- i=2855
      ("1000011100110100", "011"), -- i=2856
      ("1001011100110100", "011"), -- i=2857
      ("1010011100110100", "011"), -- i=2858
      ("1011011100110100", "011"), -- i=2859
      ("0101011100110000", "011"), -- i=2860
      ("0100011100110000", "011"), -- i=2861
      ("1000011100110101", "011"), -- i=2862
      ("1001011100110101", "011"), -- i=2863
      ("1010011100110101", "011"), -- i=2864
      ("1011011100110101", "011"), -- i=2865
      ("0101011100110000", "011"), -- i=2866
      ("0100011100110000", "011"), -- i=2867
      ("1000011100110110", "011"), -- i=2868
      ("1001011100110110", "011"), -- i=2869
      ("1010011100110110", "011"), -- i=2870
      ("1011011100110110", "011"), -- i=2871
      ("0101011100110000", "011"), -- i=2872
      ("0100011100110000", "011"), -- i=2873
      ("1000011100110111", "011"), -- i=2874
      ("1001011100110111", "011"), -- i=2875
      ("1010011100110111", "011"), -- i=2876
      ("1011011100110111", "011"), -- i=2877
      ("0101011100110000", "011"), -- i=2878
      ("0100011100110000", "011"), -- i=2879
      ("1000011101000000", "100"), -- i=2880
      ("1001011101000000", "100"), -- i=2881
      ("1010011101000000", "100"), -- i=2882
      ("1011011101000000", "100"), -- i=2883
      ("0101011101000000", "100"), -- i=2884
      ("0100011101000000", "100"), -- i=2885
      ("1000011101000001", "100"), -- i=2886
      ("1001011101000001", "100"), -- i=2887
      ("1010011101000001", "100"), -- i=2888
      ("1011011101000001", "100"), -- i=2889
      ("0101011101000000", "100"), -- i=2890
      ("0100011101000000", "100"), -- i=2891
      ("1000011101000010", "100"), -- i=2892
      ("1001011101000010", "100"), -- i=2893
      ("1010011101000010", "100"), -- i=2894
      ("1011011101000010", "100"), -- i=2895
      ("0101011101000000", "100"), -- i=2896
      ("0100011101000000", "100"), -- i=2897
      ("1000011101000011", "100"), -- i=2898
      ("1001011101000011", "100"), -- i=2899
      ("1010011101000011", "100"), -- i=2900
      ("1011011101000011", "100"), -- i=2901
      ("0101011101000000", "100"), -- i=2902
      ("0100011101000000", "100"), -- i=2903
      ("1000011101000100", "100"), -- i=2904
      ("1001011101000100", "100"), -- i=2905
      ("1010011101000100", "100"), -- i=2906
      ("1011011101000100", "100"), -- i=2907
      ("0101011101000000", "100"), -- i=2908
      ("0100011101000000", "100"), -- i=2909
      ("1000011101000101", "100"), -- i=2910
      ("1001011101000101", "100"), -- i=2911
      ("1010011101000101", "100"), -- i=2912
      ("1011011101000101", "100"), -- i=2913
      ("0101011101000000", "100"), -- i=2914
      ("0100011101000000", "100"), -- i=2915
      ("1000011101000110", "100"), -- i=2916
      ("1001011101000110", "100"), -- i=2917
      ("1010011101000110", "100"), -- i=2918
      ("1011011101000110", "100"), -- i=2919
      ("0101011101000000", "100"), -- i=2920
      ("0100011101000000", "100"), -- i=2921
      ("1000011101000111", "100"), -- i=2922
      ("1001011101000111", "100"), -- i=2923
      ("1010011101000111", "100"), -- i=2924
      ("1011011101000111", "100"), -- i=2925
      ("0101011101000000", "100"), -- i=2926
      ("0100011101000000", "100"), -- i=2927
      ("1000011101010000", "101"), -- i=2928
      ("1001011101010000", "101"), -- i=2929
      ("1010011101010000", "101"), -- i=2930
      ("1011011101010000", "101"), -- i=2931
      ("0101011101010000", "101"), -- i=2932
      ("0100011101010000", "101"), -- i=2933
      ("1000011101010001", "101"), -- i=2934
      ("1001011101010001", "101"), -- i=2935
      ("1010011101010001", "101"), -- i=2936
      ("1011011101010001", "101"), -- i=2937
      ("0101011101010000", "101"), -- i=2938
      ("0100011101010000", "101"), -- i=2939
      ("1000011101010010", "101"), -- i=2940
      ("1001011101010010", "101"), -- i=2941
      ("1010011101010010", "101"), -- i=2942
      ("1011011101010010", "101"), -- i=2943
      ("0101011101010000", "101"), -- i=2944
      ("0100011101010000", "101"), -- i=2945
      ("1000011101010011", "101"), -- i=2946
      ("1001011101010011", "101"), -- i=2947
      ("1010011101010011", "101"), -- i=2948
      ("1011011101010011", "101"), -- i=2949
      ("0101011101010000", "101"), -- i=2950
      ("0100011101010000", "101"), -- i=2951
      ("1000011101010100", "101"), -- i=2952
      ("1001011101010100", "101"), -- i=2953
      ("1010011101010100", "101"), -- i=2954
      ("1011011101010100", "101"), -- i=2955
      ("0101011101010000", "101"), -- i=2956
      ("0100011101010000", "101"), -- i=2957
      ("1000011101010101", "101"), -- i=2958
      ("1001011101010101", "101"), -- i=2959
      ("1010011101010101", "101"), -- i=2960
      ("1011011101010101", "101"), -- i=2961
      ("0101011101010000", "101"), -- i=2962
      ("0100011101010000", "101"), -- i=2963
      ("1000011101010110", "101"), -- i=2964
      ("1001011101010110", "101"), -- i=2965
      ("1010011101010110", "101"), -- i=2966
      ("1011011101010110", "101"), -- i=2967
      ("0101011101010000", "101"), -- i=2968
      ("0100011101010000", "101"), -- i=2969
      ("1000011101010111", "101"), -- i=2970
      ("1001011101010111", "101"), -- i=2971
      ("1010011101010111", "101"), -- i=2972
      ("1011011101010111", "101"), -- i=2973
      ("0101011101010000", "101"), -- i=2974
      ("0100011101010000", "101"), -- i=2975
      ("1000011101100000", "110"), -- i=2976
      ("1001011101100000", "110"), -- i=2977
      ("1010011101100000", "110"), -- i=2978
      ("1011011101100000", "110"), -- i=2979
      ("0101011101100000", "110"), -- i=2980
      ("0100011101100000", "110"), -- i=2981
      ("1000011101100001", "110"), -- i=2982
      ("1001011101100001", "110"), -- i=2983
      ("1010011101100001", "110"), -- i=2984
      ("1011011101100001", "110"), -- i=2985
      ("0101011101100000", "110"), -- i=2986
      ("0100011101100000", "110"), -- i=2987
      ("1000011101100010", "110"), -- i=2988
      ("1001011101100010", "110"), -- i=2989
      ("1010011101100010", "110"), -- i=2990
      ("1011011101100010", "110"), -- i=2991
      ("0101011101100000", "110"), -- i=2992
      ("0100011101100000", "110"), -- i=2993
      ("1000011101100011", "110"), -- i=2994
      ("1001011101100011", "110"), -- i=2995
      ("1010011101100011", "110"), -- i=2996
      ("1011011101100011", "110"), -- i=2997
      ("0101011101100000", "110"), -- i=2998
      ("0100011101100000", "110"), -- i=2999
      ("1000011101100100", "110"), -- i=3000
      ("1001011101100100", "110"), -- i=3001
      ("1010011101100100", "110"), -- i=3002
      ("1011011101100100", "110"), -- i=3003
      ("0101011101100000", "110"), -- i=3004
      ("0100011101100000", "110"), -- i=3005
      ("1000011101100101", "110"), -- i=3006
      ("1001011101100101", "110"), -- i=3007
      ("1010011101100101", "110"), -- i=3008
      ("1011011101100101", "110"), -- i=3009
      ("0101011101100000", "110"), -- i=3010
      ("0100011101100000", "110"), -- i=3011
      ("1000011101100110", "110"), -- i=3012
      ("1001011101100110", "110"), -- i=3013
      ("1010011101100110", "110"), -- i=3014
      ("1011011101100110", "110"), -- i=3015
      ("0101011101100000", "110"), -- i=3016
      ("0100011101100000", "110"), -- i=3017
      ("1000011101100111", "110"), -- i=3018
      ("1001011101100111", "110"), -- i=3019
      ("1010011101100111", "110"), -- i=3020
      ("1011011101100111", "110"), -- i=3021
      ("0101011101100000", "110"), -- i=3022
      ("0100011101100000", "110"), -- i=3023
      ("1000011101110000", "111"), -- i=3024
      ("1001011101110000", "111"), -- i=3025
      ("1010011101110000", "111"), -- i=3026
      ("1011011101110000", "111"), -- i=3027
      ("0101011101110000", "111"), -- i=3028
      ("0100011101110000", "111"), -- i=3029
      ("1000011101110001", "111"), -- i=3030
      ("1001011101110001", "111"), -- i=3031
      ("1010011101110001", "111"), -- i=3032
      ("1011011101110001", "111"), -- i=3033
      ("0101011101110000", "111"), -- i=3034
      ("0100011101110000", "111"), -- i=3035
      ("1000011101110010", "111"), -- i=3036
      ("1001011101110010", "111"), -- i=3037
      ("1010011101110010", "111"), -- i=3038
      ("1011011101110010", "111"), -- i=3039
      ("0101011101110000", "111"), -- i=3040
      ("0100011101110000", "111"), -- i=3041
      ("1000011101110011", "111"), -- i=3042
      ("1001011101110011", "111"), -- i=3043
      ("1010011101110011", "111"), -- i=3044
      ("1011011101110011", "111"), -- i=3045
      ("0101011101110000", "111"), -- i=3046
      ("0100011101110000", "111"), -- i=3047
      ("1000011101110100", "111"), -- i=3048
      ("1001011101110100", "111"), -- i=3049
      ("1010011101110100", "111"), -- i=3050
      ("1011011101110100", "111"), -- i=3051
      ("0101011101110000", "111"), -- i=3052
      ("0100011101110000", "111"), -- i=3053
      ("1000011101110101", "111"), -- i=3054
      ("1001011101110101", "111"), -- i=3055
      ("1010011101110101", "111"), -- i=3056
      ("1011011101110101", "111"), -- i=3057
      ("0101011101110000", "111"), -- i=3058
      ("0100011101110000", "111"), -- i=3059
      ("1000011101110110", "111"), -- i=3060
      ("1001011101110110", "111"), -- i=3061
      ("1010011101110110", "111"), -- i=3062
      ("1011011101110110", "111"), -- i=3063
      ("0101011101110000", "111"), -- i=3064
      ("0100011101110000", "111"), -- i=3065
      ("1000011101110111", "111"), -- i=3066
      ("1001011101110111", "111"), -- i=3067
      ("1010011101110111", "111"), -- i=3068
      ("1011011101110111", "111"), -- i=3069
      ("0101011101110000", "111"), -- i=3070
      ("0100011101110000", "111"));
  begin
    for i in patterns'range loop
      INST <= patterns(i).INST;
      wait for 10 ns;
      assert std_match(ALUOP, patterns(i).ALUOP) OR (ALUOP = "ZZ" AND patterns(i).ALUOP = "ZZ")
        report "wrong value for ALUOP, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).ALUOP) & ", found " & to_string(ALUOP) severity error;assert std_match(RS1, patterns(i).RS1) OR (RS1 = "ZZZ" AND patterns(i).RS1 = "ZZZ")
        report "wrong value for RS1, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).RS1) & ", found " & to_string(RS1) severity error;assert std_match(RS2, patterns(i).RS2) OR (RS2 = "ZZZ" AND patterns(i).RS2 = "ZZZ")
        report "wrong value for RS2, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).RS2) & ", found " & to_string(RS2) severity error;assert std_match(WS, patterns(i).WS) OR (WS = "ZZZ" AND patterns(i).WS = "ZZZ")
        report "wrong value for WS, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).WS) & ", found " & to_string(WS) severity error;assert std_match(STR, patterns(i).STR) OR (STR = 'Z' AND patterns(i).STR = 'Z')
        report "wrong value for STR, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).STR) & ", found " & std_logic'image(STR) severity error;assert std_match(WE, patterns(i).WE) OR (WE = 'Z' AND patterns(i).WE = 'Z')
        report "wrong value for WE, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).WE) & ", found " & std_logic'image(WE) severity error;assert std_match(DMUX, patterns(i).DMUX) OR (DMUX = "ZZ" AND patterns(i).DMUX = "ZZ")
        report "wrong value for DMUX, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).DMUX) & ", found " & to_string(DMUX) severity error;assert std_match(LDR, patterns(i).LDR) OR (LDR = 'Z' AND patterns(i).LDR = 'Z')
        report "wrong value for LDR, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).LDR) & ", found " & std_logic'image(LDR) severity error;end loop;
    wait;
  end process;
end behav;
