--  A testbench for control_unit_LDR_tb
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity control_unit_LDR_tb is
end control_unit_LDR_tb;

architecture behav of control_unit_LDR_tb is
  component main
    port (
      INST: in std_logic_vector(15 downto 0);
      ALUOP: out std_logic_vector(1 downto 0);
      RS1: out std_logic_vector(2 downto 0);
      RS2: out std_logic_vector(2 downto 0);
      WS: out std_logic_vector(2 downto 0);
      STR: out std_logic;
      WE: out std_logic;
      DMUX: out std_logic_vector(1 downto 0);
      LDR: out std_logic);
  end component;

  signal INST : std_logic_vector(15 downto 0);
  signal ALUOP : std_logic_vector(1 downto 0);
  signal RS1 : std_logic_vector(2 downto 0);
  signal RS2 : std_logic_vector(2 downto 0);
  signal WS : std_logic_vector(2 downto 0);
  signal STR : std_logic;
  signal WE : std_logic;
  signal DMUX : std_logic_vector(1 downto 0);
  signal LDR : std_logic;
  function to_string ( a: std_logic_vector) return string is
      variable b : string (1 to a'length) := (others => NUL);
      variable stri : integer := 1; 
  begin
      for i in a'range loop
          b(stri) := std_logic'image(a((i)))(2);
      stri := stri+1;
      end loop;
      return b;
  end function;
begin
  main_0 : main port map (
    INST => INST,
    ALUOP => ALUOP,
    RS1 => RS1,
    RS2 => RS2,
    WS => WS,
    STR => STR,
    WE => WE,
    DMUX => DMUX,
    LDR => LDR );
  process
    type pattern_type is record
      INST : std_logic_vector(15 downto 0);
      LDR : std_logic;
    end record;
    type pattern_array is array (natural range <>) of pattern_type;
    constant patterns : pattern_array := (
      ("1000000000000000", '-'), -- i=0
      ("1001000000000000", '-'), -- i=1
      ("1010000000000000", '-'), -- i=2
      ("1011000000000000", '-'), -- i=3
      ("0101000000000000", '1'), -- i=4
      ("0100000000000000", '-'), -- i=5
      ("0000000001000010", '-'), -- i=6
      ("1000000000000001", '-'), -- i=7
      ("1001000000000001", '-'), -- i=8
      ("1010000000000001", '-'), -- i=9
      ("1011000000000001", '-'), -- i=10
      ("0101000000000000", '1'), -- i=11
      ("0100000000000000", '-'), -- i=12
      ("0000000010011010", '-'), -- i=13
      ("1000000000000010", '-'), -- i=14
      ("1001000000000010", '-'), -- i=15
      ("1010000000000010", '-'), -- i=16
      ("1011000000000010", '-'), -- i=17
      ("0101000000000000", '1'), -- i=18
      ("0100000000000000", '-'), -- i=19
      ("0000000000101100", '-'), -- i=20
      ("1000000000000011", '-'), -- i=21
      ("1001000000000011", '-'), -- i=22
      ("1010000000000011", '-'), -- i=23
      ("1011000000000011", '-'), -- i=24
      ("0101000000000000", '1'), -- i=25
      ("0100000000000000", '-'), -- i=26
      ("0000000001001011", '-'), -- i=27
      ("1000000000000100", '-'), -- i=28
      ("1001000000000100", '-'), -- i=29
      ("1010000000000100", '-'), -- i=30
      ("1011000000000100", '-'), -- i=31
      ("0101000000000000", '1'), -- i=32
      ("0100000000000000", '-'), -- i=33
      ("0000000011101110", '-'), -- i=34
      ("1000000000000101", '-'), -- i=35
      ("1001000000000101", '-'), -- i=36
      ("1010000000000101", '-'), -- i=37
      ("1011000000000101", '-'), -- i=38
      ("0101000000000000", '1'), -- i=39
      ("0100000000000000", '-'), -- i=40
      ("0000000001101001", '-'), -- i=41
      ("1000000000000110", '-'), -- i=42
      ("1001000000000110", '-'), -- i=43
      ("1010000000000110", '-'), -- i=44
      ("1011000000000110", '-'), -- i=45
      ("0101000000000000", '1'), -- i=46
      ("0100000000000000", '-'), -- i=47
      ("0000000001011011", '-'), -- i=48
      ("1000000000000111", '-'), -- i=49
      ("1001000000000111", '-'), -- i=50
      ("1010000000000111", '-'), -- i=51
      ("1011000000000111", '-'), -- i=52
      ("0101000000000000", '1'), -- i=53
      ("0100000000000000", '-'), -- i=54
      ("0000000000100011", '-'), -- i=55
      ("1000000000010000", '-'), -- i=56
      ("1001000000010000", '-'), -- i=57
      ("1010000000010000", '-'), -- i=58
      ("1011000000010000", '-'), -- i=59
      ("0101000000010000", '1'), -- i=60
      ("0100000000010000", '-'), -- i=61
      ("0000000010111111", '-'), -- i=62
      ("1000000000010001", '-'), -- i=63
      ("1001000000010001", '-'), -- i=64
      ("1010000000010001", '-'), -- i=65
      ("1011000000010001", '-'), -- i=66
      ("0101000000010000", '1'), -- i=67
      ("0100000000010000", '-'), -- i=68
      ("0000000010000111", '-'), -- i=69
      ("1000000000010010", '-'), -- i=70
      ("1001000000010010", '-'), -- i=71
      ("1010000000010010", '-'), -- i=72
      ("1011000000010010", '-'), -- i=73
      ("0101000000010000", '1'), -- i=74
      ("0100000000010000", '-'), -- i=75
      ("0000000000101101", '-'), -- i=76
      ("1000000000010011", '-'), -- i=77
      ("1001000000010011", '-'), -- i=78
      ("1010000000010011", '-'), -- i=79
      ("1011000000010011", '-'), -- i=80
      ("0101000000010000", '1'), -- i=81
      ("0100000000010000", '-'), -- i=82
      ("0000000001101110", '-'), -- i=83
      ("1000000000010100", '-'), -- i=84
      ("1001000000010100", '-'), -- i=85
      ("1010000000010100", '-'), -- i=86
      ("1011000000010100", '-'), -- i=87
      ("0101000000010000", '1'), -- i=88
      ("0100000000010000", '-'), -- i=89
      ("0000000010010101", '-'), -- i=90
      ("1000000000010101", '-'), -- i=91
      ("1001000000010101", '-'), -- i=92
      ("1010000000010101", '-'), -- i=93
      ("1011000000010101", '-'), -- i=94
      ("0101000000010000", '1'), -- i=95
      ("0100000000010000", '-'), -- i=96
      ("0000000000100100", '-'), -- i=97
      ("1000000000010110", '-'), -- i=98
      ("1001000000010110", '-'), -- i=99
      ("1010000000010110", '-'), -- i=100
      ("1011000000010110", '-'), -- i=101
      ("0101000000010000", '1'), -- i=102
      ("0100000000010000", '-'), -- i=103
      ("0000000000111011", '-'), -- i=104
      ("1000000000010111", '-'), -- i=105
      ("1001000000010111", '-'), -- i=106
      ("1010000000010111", '-'), -- i=107
      ("1011000000010111", '-'), -- i=108
      ("0101000000010000", '1'), -- i=109
      ("0100000000010000", '-'), -- i=110
      ("0000000001111111", '-'), -- i=111
      ("1000000000100000", '-'), -- i=112
      ("1001000000100000", '-'), -- i=113
      ("1010000000100000", '-'), -- i=114
      ("1011000000100000", '-'), -- i=115
      ("0101000000100000", '1'), -- i=116
      ("0100000000100000", '-'), -- i=117
      ("0000000000111011", '-'), -- i=118
      ("1000000000100001", '-'), -- i=119
      ("1001000000100001", '-'), -- i=120
      ("1010000000100001", '-'), -- i=121
      ("1011000000100001", '-'), -- i=122
      ("0101000000100000", '1'), -- i=123
      ("0100000000100000", '-'), -- i=124
      ("0000000011010101", '-'), -- i=125
      ("1000000000100010", '-'), -- i=126
      ("1001000000100010", '-'), -- i=127
      ("1010000000100010", '-'), -- i=128
      ("1011000000100010", '-'), -- i=129
      ("0101000000100000", '1'), -- i=130
      ("0100000000100000", '-'), -- i=131
      ("0000000001110110", '-'), -- i=132
      ("1000000000100011", '-'), -- i=133
      ("1001000000100011", '-'), -- i=134
      ("1010000000100011", '-'), -- i=135
      ("1011000000100011", '-'), -- i=136
      ("0101000000100000", '1'), -- i=137
      ("0100000000100000", '-'), -- i=138
      ("0000000000111010", '-'), -- i=139
      ("1000000000100100", '-'), -- i=140
      ("1001000000100100", '-'), -- i=141
      ("1010000000100100", '-'), -- i=142
      ("1011000000100100", '-'), -- i=143
      ("0101000000100000", '1'), -- i=144
      ("0100000000100000", '-'), -- i=145
      ("0000000010000100", '-'), -- i=146
      ("1000000000100101", '-'), -- i=147
      ("1001000000100101", '-'), -- i=148
      ("1010000000100101", '-'), -- i=149
      ("1011000000100101", '-'), -- i=150
      ("0101000000100000", '1'), -- i=151
      ("0100000000100000", '-'), -- i=152
      ("0000000001010011", '-'), -- i=153
      ("1000000000100110", '-'), -- i=154
      ("1001000000100110", '-'), -- i=155
      ("1010000000100110", '-'), -- i=156
      ("1011000000100110", '-'), -- i=157
      ("0101000000100000", '1'), -- i=158
      ("0100000000100000", '-'), -- i=159
      ("0000000011000101", '-'), -- i=160
      ("1000000000100111", '-'), -- i=161
      ("1001000000100111", '-'), -- i=162
      ("1010000000100111", '-'), -- i=163
      ("1011000000100111", '-'), -- i=164
      ("0101000000100000", '1'), -- i=165
      ("0100000000100000", '-'), -- i=166
      ("0000000001110000", '-'), -- i=167
      ("1000000000110000", '-'), -- i=168
      ("1001000000110000", '-'), -- i=169
      ("1010000000110000", '-'), -- i=170
      ("1011000000110000", '-'), -- i=171
      ("0101000000110000", '1'), -- i=172
      ("0100000000110000", '-'), -- i=173
      ("0000000000110010", '-'), -- i=174
      ("1000000000110001", '-'), -- i=175
      ("1001000000110001", '-'), -- i=176
      ("1010000000110001", '-'), -- i=177
      ("1011000000110001", '-'), -- i=178
      ("0101000000110000", '1'), -- i=179
      ("0100000000110000", '-'), -- i=180
      ("0000000001101011", '-'), -- i=181
      ("1000000000110010", '-'), -- i=182
      ("1001000000110010", '-'), -- i=183
      ("1010000000110010", '-'), -- i=184
      ("1011000000110010", '-'), -- i=185
      ("0101000000110000", '1'), -- i=186
      ("0100000000110000", '-'), -- i=187
      ("0000000010001010", '-'), -- i=188
      ("1000000000110011", '-'), -- i=189
      ("1001000000110011", '-'), -- i=190
      ("1010000000110011", '-'), -- i=191
      ("1011000000110011", '-'), -- i=192
      ("0101000000110000", '1'), -- i=193
      ("0100000000110000", '-'), -- i=194
      ("0000000000100111", '-'), -- i=195
      ("1000000000110100", '-'), -- i=196
      ("1001000000110100", '-'), -- i=197
      ("1010000000110100", '-'), -- i=198
      ("1011000000110100", '-'), -- i=199
      ("0101000000110000", '1'), -- i=200
      ("0100000000110000", '-'), -- i=201
      ("0000000000111000", '-'), -- i=202
      ("1000000000110101", '-'), -- i=203
      ("1001000000110101", '-'), -- i=204
      ("1010000000110101", '-'), -- i=205
      ("1011000000110101", '-'), -- i=206
      ("0101000000110000", '1'), -- i=207
      ("0100000000110000", '-'), -- i=208
      ("0000000001000001", '-'), -- i=209
      ("1000000000110110", '-'), -- i=210
      ("1001000000110110", '-'), -- i=211
      ("1010000000110110", '-'), -- i=212
      ("1011000000110110", '-'), -- i=213
      ("0101000000110000", '1'), -- i=214
      ("0100000000110000", '-'), -- i=215
      ("0000000010100100", '-'), -- i=216
      ("1000000000110111", '-'), -- i=217
      ("1001000000110111", '-'), -- i=218
      ("1010000000110111", '-'), -- i=219
      ("1011000000110111", '-'), -- i=220
      ("0101000000110000", '1'), -- i=221
      ("0100000000110000", '-'), -- i=222
      ("0000000010011011", '-'), -- i=223
      ("1000000001000000", '-'), -- i=224
      ("1001000001000000", '-'), -- i=225
      ("1010000001000000", '-'), -- i=226
      ("1011000001000000", '-'), -- i=227
      ("0101000001000000", '1'), -- i=228
      ("0100000001000000", '-'), -- i=229
      ("0000000011110000", '-'), -- i=230
      ("1000000001000001", '-'), -- i=231
      ("1001000001000001", '-'), -- i=232
      ("1010000001000001", '-'), -- i=233
      ("1011000001000001", '-'), -- i=234
      ("0101000001000000", '1'), -- i=235
      ("0100000001000000", '-'), -- i=236
      ("0000000000001011", '-'), -- i=237
      ("1000000001000010", '-'), -- i=238
      ("1001000001000010", '-'), -- i=239
      ("1010000001000010", '-'), -- i=240
      ("1011000001000010", '-'), -- i=241
      ("0101000001000000", '1'), -- i=242
      ("0100000001000000", '-'), -- i=243
      ("0000000010000111", '-'), -- i=244
      ("1000000001000011", '-'), -- i=245
      ("1001000001000011", '-'), -- i=246
      ("1010000001000011", '-'), -- i=247
      ("1011000001000011", '-'), -- i=248
      ("0101000001000000", '1'), -- i=249
      ("0100000001000000", '-'), -- i=250
      ("0000000001011000", '-'), -- i=251
      ("1000000001000100", '-'), -- i=252
      ("1001000001000100", '-'), -- i=253
      ("1010000001000100", '-'), -- i=254
      ("1011000001000100", '-'), -- i=255
      ("0101000001000000", '1'), -- i=256
      ("0100000001000000", '-'), -- i=257
      ("0000000000111111", '-'), -- i=258
      ("1000000001000101", '-'), -- i=259
      ("1001000001000101", '-'), -- i=260
      ("1010000001000101", '-'), -- i=261
      ("1011000001000101", '-'), -- i=262
      ("0101000001000000", '1'), -- i=263
      ("0100000001000000", '-'), -- i=264
      ("0000000000010100", '-'), -- i=265
      ("1000000001000110", '-'), -- i=266
      ("1001000001000110", '-'), -- i=267
      ("1010000001000110", '-'), -- i=268
      ("1011000001000110", '-'), -- i=269
      ("0101000001000000", '1'), -- i=270
      ("0100000001000000", '-'), -- i=271
      ("0000000000110111", '-'), -- i=272
      ("1000000001000111", '-'), -- i=273
      ("1001000001000111", '-'), -- i=274
      ("1010000001000111", '-'), -- i=275
      ("1011000001000111", '-'), -- i=276
      ("0101000001000000", '1'), -- i=277
      ("0100000001000000", '-'), -- i=278
      ("0000000011110001", '-'), -- i=279
      ("1000000001010000", '-'), -- i=280
      ("1001000001010000", '-'), -- i=281
      ("1010000001010000", '-'), -- i=282
      ("1011000001010000", '-'), -- i=283
      ("0101000001010000", '1'), -- i=284
      ("0100000001010000", '-'), -- i=285
      ("0000000010011001", '-'), -- i=286
      ("1000000001010001", '-'), -- i=287
      ("1001000001010001", '-'), -- i=288
      ("1010000001010001", '-'), -- i=289
      ("1011000001010001", '-'), -- i=290
      ("0101000001010000", '1'), -- i=291
      ("0100000001010000", '-'), -- i=292
      ("0000000001100110", '-'), -- i=293
      ("1000000001010010", '-'), -- i=294
      ("1001000001010010", '-'), -- i=295
      ("1010000001010010", '-'), -- i=296
      ("1011000001010010", '-'), -- i=297
      ("0101000001010000", '1'), -- i=298
      ("0100000001010000", '-'), -- i=299
      ("0000000011011010", '-'), -- i=300
      ("1000000001010011", '-'), -- i=301
      ("1001000001010011", '-'), -- i=302
      ("1010000001010011", '-'), -- i=303
      ("1011000001010011", '-'), -- i=304
      ("0101000001010000", '1'), -- i=305
      ("0100000001010000", '-'), -- i=306
      ("0000000011110000", '-'), -- i=307
      ("1000000001010100", '-'), -- i=308
      ("1001000001010100", '-'), -- i=309
      ("1010000001010100", '-'), -- i=310
      ("1011000001010100", '-'), -- i=311
      ("0101000001010000", '1'), -- i=312
      ("0100000001010000", '-'), -- i=313
      ("0000000001010100", '-'), -- i=314
      ("1000000001010101", '-'), -- i=315
      ("1001000001010101", '-'), -- i=316
      ("1010000001010101", '-'), -- i=317
      ("1011000001010101", '-'), -- i=318
      ("0101000001010000", '1'), -- i=319
      ("0100000001010000", '-'), -- i=320
      ("0000000010110000", '-'), -- i=321
      ("1000000001010110", '-'), -- i=322
      ("1001000001010110", '-'), -- i=323
      ("1010000001010110", '-'), -- i=324
      ("1011000001010110", '-'), -- i=325
      ("0101000001010000", '1'), -- i=326
      ("0100000001010000", '-'), -- i=327
      ("0000000011101110", '-'), -- i=328
      ("1000000001010111", '-'), -- i=329
      ("1001000001010111", '-'), -- i=330
      ("1010000001010111", '-'), -- i=331
      ("1011000001010111", '-'), -- i=332
      ("0101000001010000", '1'), -- i=333
      ("0100000001010000", '-'), -- i=334
      ("0000000001001011", '-'), -- i=335
      ("1000000001100000", '-'), -- i=336
      ("1001000001100000", '-'), -- i=337
      ("1010000001100000", '-'), -- i=338
      ("1011000001100000", '-'), -- i=339
      ("0101000001100000", '1'), -- i=340
      ("0100000001100000", '-'), -- i=341
      ("0000000011000000", '-'), -- i=342
      ("1000000001100001", '-'), -- i=343
      ("1001000001100001", '-'), -- i=344
      ("1010000001100001", '-'), -- i=345
      ("1011000001100001", '-'), -- i=346
      ("0101000001100000", '1'), -- i=347
      ("0100000001100000", '-'), -- i=348
      ("0000000000100110", '-'), -- i=349
      ("1000000001100010", '-'), -- i=350
      ("1001000001100010", '-'), -- i=351
      ("1010000001100010", '-'), -- i=352
      ("1011000001100010", '-'), -- i=353
      ("0101000001100000", '1'), -- i=354
      ("0100000001100000", '-'), -- i=355
      ("0000000000101010", '-'), -- i=356
      ("1000000001100011", '-'), -- i=357
      ("1001000001100011", '-'), -- i=358
      ("1010000001100011", '-'), -- i=359
      ("1011000001100011", '-'), -- i=360
      ("0101000001100000", '1'), -- i=361
      ("0100000001100000", '-'), -- i=362
      ("0000000001101101", '-'), -- i=363
      ("1000000001100100", '-'), -- i=364
      ("1001000001100100", '-'), -- i=365
      ("1010000001100100", '-'), -- i=366
      ("1011000001100100", '-'), -- i=367
      ("0101000001100000", '1'), -- i=368
      ("0100000001100000", '-'), -- i=369
      ("0000000000001010", '-'), -- i=370
      ("1000000001100101", '-'), -- i=371
      ("1001000001100101", '-'), -- i=372
      ("1010000001100101", '-'), -- i=373
      ("1011000001100101", '-'), -- i=374
      ("0101000001100000", '1'), -- i=375
      ("0100000001100000", '-'), -- i=376
      ("0000000011010001", '-'), -- i=377
      ("1000000001100110", '-'), -- i=378
      ("1001000001100110", '-'), -- i=379
      ("1010000001100110", '-'), -- i=380
      ("1011000001100110", '-'), -- i=381
      ("0101000001100000", '1'), -- i=382
      ("0100000001100000", '-'), -- i=383
      ("0000000001100111", '-'), -- i=384
      ("1000000001100111", '-'), -- i=385
      ("1001000001100111", '-'), -- i=386
      ("1010000001100111", '-'), -- i=387
      ("1011000001100111", '-'), -- i=388
      ("0101000001100000", '1'), -- i=389
      ("0100000001100000", '-'), -- i=390
      ("0000000000000000", '-'), -- i=391
      ("1000000001110000", '-'), -- i=392
      ("1001000001110000", '-'), -- i=393
      ("1010000001110000", '-'), -- i=394
      ("1011000001110000", '-'), -- i=395
      ("0101000001110000", '1'), -- i=396
      ("0100000001110000", '-'), -- i=397
      ("0000000000001011", '-'), -- i=398
      ("1000000001110001", '-'), -- i=399
      ("1001000001110001", '-'), -- i=400
      ("1010000001110001", '-'), -- i=401
      ("1011000001110001", '-'), -- i=402
      ("0101000001110000", '1'), -- i=403
      ("0100000001110000", '-'), -- i=404
      ("0000000010000010", '-'), -- i=405
      ("1000000001110010", '-'), -- i=406
      ("1001000001110010", '-'), -- i=407
      ("1010000001110010", '-'), -- i=408
      ("1011000001110010", '-'), -- i=409
      ("0101000001110000", '1'), -- i=410
      ("0100000001110000", '-'), -- i=411
      ("0000000000010110", '-'), -- i=412
      ("1000000001110011", '-'), -- i=413
      ("1001000001110011", '-'), -- i=414
      ("1010000001110011", '-'), -- i=415
      ("1011000001110011", '-'), -- i=416
      ("0101000001110000", '1'), -- i=417
      ("0100000001110000", '-'), -- i=418
      ("0000000000001001", '-'), -- i=419
      ("1000000001110100", '-'), -- i=420
      ("1001000001110100", '-'), -- i=421
      ("1010000001110100", '-'), -- i=422
      ("1011000001110100", '-'), -- i=423
      ("0101000001110000", '1'), -- i=424
      ("0100000001110000", '-'), -- i=425
      ("0000000010101011", '-'), -- i=426
      ("1000000001110101", '-'), -- i=427
      ("1001000001110101", '-'), -- i=428
      ("1010000001110101", '-'), -- i=429
      ("1011000001110101", '-'), -- i=430
      ("0101000001110000", '1'), -- i=431
      ("0100000001110000", '-'), -- i=432
      ("0000000011111010", '-'), -- i=433
      ("1000000001110110", '-'), -- i=434
      ("1001000001110110", '-'), -- i=435
      ("1010000001110110", '-'), -- i=436
      ("1011000001110110", '-'), -- i=437
      ("0101000001110000", '1'), -- i=438
      ("0100000001110000", '-'), -- i=439
      ("0000000000000111", '-'), -- i=440
      ("1000000001110111", '-'), -- i=441
      ("1001000001110111", '-'), -- i=442
      ("1010000001110111", '-'), -- i=443
      ("1011000001110111", '-'), -- i=444
      ("0101000001110000", '1'), -- i=445
      ("0100000001110000", '-'), -- i=446
      ("0000000010011111", '-'), -- i=447
      ("1000000100000000", '-'), -- i=448
      ("1001000100000000", '-'), -- i=449
      ("1010000100000000", '-'), -- i=450
      ("1011000100000000", '-'), -- i=451
      ("0101000100000000", '1'), -- i=452
      ("0100000100000000", '-'), -- i=453
      ("0000000111001010", '-'), -- i=454
      ("1000000100000001", '-'), -- i=455
      ("1001000100000001", '-'), -- i=456
      ("1010000100000001", '-'), -- i=457
      ("1011000100000001", '-'), -- i=458
      ("0101000100000000", '1'), -- i=459
      ("0100000100000000", '-'), -- i=460
      ("0000000111111100", '-'), -- i=461
      ("1000000100000010", '-'), -- i=462
      ("1001000100000010", '-'), -- i=463
      ("1010000100000010", '-'), -- i=464
      ("1011000100000010", '-'), -- i=465
      ("0101000100000000", '1'), -- i=466
      ("0100000100000000", '-'), -- i=467
      ("0000000110101001", '-'), -- i=468
      ("1000000100000011", '-'), -- i=469
      ("1001000100000011", '-'), -- i=470
      ("1010000100000011", '-'), -- i=471
      ("1011000100000011", '-'), -- i=472
      ("0101000100000000", '1'), -- i=473
      ("0100000100000000", '-'), -- i=474
      ("0000000101100000", '-'), -- i=475
      ("1000000100000100", '-'), -- i=476
      ("1001000100000100", '-'), -- i=477
      ("1010000100000100", '-'), -- i=478
      ("1011000100000100", '-'), -- i=479
      ("0101000100000000", '1'), -- i=480
      ("0100000100000000", '-'), -- i=481
      ("0000000100111000", '-'), -- i=482
      ("1000000100000101", '-'), -- i=483
      ("1001000100000101", '-'), -- i=484
      ("1010000100000101", '-'), -- i=485
      ("1011000100000101", '-'), -- i=486
      ("0101000100000000", '1'), -- i=487
      ("0100000100000000", '-'), -- i=488
      ("0000000100001101", '-'), -- i=489
      ("1000000100000110", '-'), -- i=490
      ("1001000100000110", '-'), -- i=491
      ("1010000100000110", '-'), -- i=492
      ("1011000100000110", '-'), -- i=493
      ("0101000100000000", '1'), -- i=494
      ("0100000100000000", '-'), -- i=495
      ("0000000100010001", '-'), -- i=496
      ("1000000100000111", '-'), -- i=497
      ("1001000100000111", '-'), -- i=498
      ("1010000100000111", '-'), -- i=499
      ("1011000100000111", '-'), -- i=500
      ("0101000100000000", '1'), -- i=501
      ("0100000100000000", '-'), -- i=502
      ("0000000100101010", '-'), -- i=503
      ("1000000100010000", '-'), -- i=504
      ("1001000100010000", '-'), -- i=505
      ("1010000100010000", '-'), -- i=506
      ("1011000100010000", '-'), -- i=507
      ("0101000100010000", '1'), -- i=508
      ("0100000100010000", '-'), -- i=509
      ("0000000101110111", '-'), -- i=510
      ("1000000100010001", '-'), -- i=511
      ("1001000100010001", '-'), -- i=512
      ("1010000100010001", '-'), -- i=513
      ("1011000100010001", '-'), -- i=514
      ("0101000100010000", '1'), -- i=515
      ("0100000100010000", '-'), -- i=516
      ("0000000101010111", '-'), -- i=517
      ("1000000100010010", '-'), -- i=518
      ("1001000100010010", '-'), -- i=519
      ("1010000100010010", '-'), -- i=520
      ("1011000100010010", '-'), -- i=521
      ("0101000100010000", '1'), -- i=522
      ("0100000100010000", '-'), -- i=523
      ("0000000110100110", '-'), -- i=524
      ("1000000100010011", '-'), -- i=525
      ("1001000100010011", '-'), -- i=526
      ("1010000100010011", '-'), -- i=527
      ("1011000100010011", '-'), -- i=528
      ("0101000100010000", '1'), -- i=529
      ("0100000100010000", '-'), -- i=530
      ("0000000111110100", '-'), -- i=531
      ("1000000100010100", '-'), -- i=532
      ("1001000100010100", '-'), -- i=533
      ("1010000100010100", '-'), -- i=534
      ("1011000100010100", '-'), -- i=535
      ("0101000100010000", '1'), -- i=536
      ("0100000100010000", '-'), -- i=537
      ("0000000111010000", '-'), -- i=538
      ("1000000100010101", '-'), -- i=539
      ("1001000100010101", '-'), -- i=540
      ("1010000100010101", '-'), -- i=541
      ("1011000100010101", '-'), -- i=542
      ("0101000100010000", '1'), -- i=543
      ("0100000100010000", '-'), -- i=544
      ("0000000110101001", '-'), -- i=545
      ("1000000100010110", '-'), -- i=546
      ("1001000100010110", '-'), -- i=547
      ("1010000100010110", '-'), -- i=548
      ("1011000100010110", '-'), -- i=549
      ("0101000100010000", '1'), -- i=550
      ("0100000100010000", '-'), -- i=551
      ("0000000101111100", '-'), -- i=552
      ("1000000100010111", '-'), -- i=553
      ("1001000100010111", '-'), -- i=554
      ("1010000100010111", '-'), -- i=555
      ("1011000100010111", '-'), -- i=556
      ("0101000100010000", '1'), -- i=557
      ("0100000100010000", '-'), -- i=558
      ("0000000110010110", '-'), -- i=559
      ("1000000100100000", '-'), -- i=560
      ("1001000100100000", '-'), -- i=561
      ("1010000100100000", '-'), -- i=562
      ("1011000100100000", '-'), -- i=563
      ("0101000100100000", '1'), -- i=564
      ("0100000100100000", '-'), -- i=565
      ("0000000110001100", '-'), -- i=566
      ("1000000100100001", '-'), -- i=567
      ("1001000100100001", '-'), -- i=568
      ("1010000100100001", '-'), -- i=569
      ("1011000100100001", '-'), -- i=570
      ("0101000100100000", '1'), -- i=571
      ("0100000100100000", '-'), -- i=572
      ("0000000111110001", '-'), -- i=573
      ("1000000100100010", '-'), -- i=574
      ("1001000100100010", '-'), -- i=575
      ("1010000100100010", '-'), -- i=576
      ("1011000100100010", '-'), -- i=577
      ("0101000100100000", '1'), -- i=578
      ("0100000100100000", '-'), -- i=579
      ("0000000100000101", '-'), -- i=580
      ("1000000100100011", '-'), -- i=581
      ("1001000100100011", '-'), -- i=582
      ("1010000100100011", '-'), -- i=583
      ("1011000100100011", '-'), -- i=584
      ("0101000100100000", '1'), -- i=585
      ("0100000100100000", '-'), -- i=586
      ("0000000101010010", '-'), -- i=587
      ("1000000100100100", '-'), -- i=588
      ("1001000100100100", '-'), -- i=589
      ("1010000100100100", '-'), -- i=590
      ("1011000100100100", '-'), -- i=591
      ("0101000100100000", '1'), -- i=592
      ("0100000100100000", '-'), -- i=593
      ("0000000111010010", '-'), -- i=594
      ("1000000100100101", '-'), -- i=595
      ("1001000100100101", '-'), -- i=596
      ("1010000100100101", '-'), -- i=597
      ("1011000100100101", '-'), -- i=598
      ("0101000100100000", '1'), -- i=599
      ("0100000100100000", '-'), -- i=600
      ("0000000110011001", '-'), -- i=601
      ("1000000100100110", '-'), -- i=602
      ("1001000100100110", '-'), -- i=603
      ("1010000100100110", '-'), -- i=604
      ("1011000100100110", '-'), -- i=605
      ("0101000100100000", '1'), -- i=606
      ("0100000100100000", '-'), -- i=607
      ("0000000100000110", '-'), -- i=608
      ("1000000100100111", '-'), -- i=609
      ("1001000100100111", '-'), -- i=610
      ("1010000100100111", '-'), -- i=611
      ("1011000100100111", '-'), -- i=612
      ("0101000100100000", '1'), -- i=613
      ("0100000100100000", '-'), -- i=614
      ("0000000101010000", '-'), -- i=615
      ("1000000100110000", '-'), -- i=616
      ("1001000100110000", '-'), -- i=617
      ("1010000100110000", '-'), -- i=618
      ("1011000100110000", '-'), -- i=619
      ("0101000100110000", '1'), -- i=620
      ("0100000100110000", '-'), -- i=621
      ("0000000100101110", '-'), -- i=622
      ("1000000100110001", '-'), -- i=623
      ("1001000100110001", '-'), -- i=624
      ("1010000100110001", '-'), -- i=625
      ("1011000100110001", '-'), -- i=626
      ("0101000100110000", '1'), -- i=627
      ("0100000100110000", '-'), -- i=628
      ("0000000111111100", '-'), -- i=629
      ("1000000100110010", '-'), -- i=630
      ("1001000100110010", '-'), -- i=631
      ("1010000100110010", '-'), -- i=632
      ("1011000100110010", '-'), -- i=633
      ("0101000100110000", '1'), -- i=634
      ("0100000100110000", '-'), -- i=635
      ("0000000101010011", '-'), -- i=636
      ("1000000100110011", '-'), -- i=637
      ("1001000100110011", '-'), -- i=638
      ("1010000100110011", '-'), -- i=639
      ("1011000100110011", '-'), -- i=640
      ("0101000100110000", '1'), -- i=641
      ("0100000100110000", '-'), -- i=642
      ("0000000111011001", '-'), -- i=643
      ("1000000100110100", '-'), -- i=644
      ("1001000100110100", '-'), -- i=645
      ("1010000100110100", '-'), -- i=646
      ("1011000100110100", '-'), -- i=647
      ("0101000100110000", '1'), -- i=648
      ("0100000100110000", '-'), -- i=649
      ("0000000110000000", '-'), -- i=650
      ("1000000100110101", '-'), -- i=651
      ("1001000100110101", '-'), -- i=652
      ("1010000100110101", '-'), -- i=653
      ("1011000100110101", '-'), -- i=654
      ("0101000100110000", '1'), -- i=655
      ("0100000100110000", '-'), -- i=656
      ("0000000100001001", '-'), -- i=657
      ("1000000100110110", '-'), -- i=658
      ("1001000100110110", '-'), -- i=659
      ("1010000100110110", '-'), -- i=660
      ("1011000100110110", '-'), -- i=661
      ("0101000100110000", '1'), -- i=662
      ("0100000100110000", '-'), -- i=663
      ("0000000101010001", '-'), -- i=664
      ("1000000100110111", '-'), -- i=665
      ("1001000100110111", '-'), -- i=666
      ("1010000100110111", '-'), -- i=667
      ("1011000100110111", '-'), -- i=668
      ("0101000100110000", '1'), -- i=669
      ("0100000100110000", '-'), -- i=670
      ("0000000100011111", '-'), -- i=671
      ("1000000101000000", '-'), -- i=672
      ("1001000101000000", '-'), -- i=673
      ("1010000101000000", '-'), -- i=674
      ("1011000101000000", '-'), -- i=675
      ("0101000101000000", '1'), -- i=676
      ("0100000101000000", '-'), -- i=677
      ("0000000110000010", '-'), -- i=678
      ("1000000101000001", '-'), -- i=679
      ("1001000101000001", '-'), -- i=680
      ("1010000101000001", '-'), -- i=681
      ("1011000101000001", '-'), -- i=682
      ("0101000101000000", '1'), -- i=683
      ("0100000101000000", '-'), -- i=684
      ("0000000101010011", '-'), -- i=685
      ("1000000101000010", '-'), -- i=686
      ("1001000101000010", '-'), -- i=687
      ("1010000101000010", '-'), -- i=688
      ("1011000101000010", '-'), -- i=689
      ("0101000101000000", '1'), -- i=690
      ("0100000101000000", '-'), -- i=691
      ("0000000111000001", '-'), -- i=692
      ("1000000101000011", '-'), -- i=693
      ("1001000101000011", '-'), -- i=694
      ("1010000101000011", '-'), -- i=695
      ("1011000101000011", '-'), -- i=696
      ("0101000101000000", '1'), -- i=697
      ("0100000101000000", '-'), -- i=698
      ("0000000101111101", '-'), -- i=699
      ("1000000101000100", '-'), -- i=700
      ("1001000101000100", '-'), -- i=701
      ("1010000101000100", '-'), -- i=702
      ("1011000101000100", '-'), -- i=703
      ("0101000101000000", '1'), -- i=704
      ("0100000101000000", '-'), -- i=705
      ("0000000100010000", '-'), -- i=706
      ("1000000101000101", '-'), -- i=707
      ("1001000101000101", '-'), -- i=708
      ("1010000101000101", '-'), -- i=709
      ("1011000101000101", '-'), -- i=710
      ("0101000101000000", '1'), -- i=711
      ("0100000101000000", '-'), -- i=712
      ("0000000100111111", '-'), -- i=713
      ("1000000101000110", '-'), -- i=714
      ("1001000101000110", '-'), -- i=715
      ("1010000101000110", '-'), -- i=716
      ("1011000101000110", '-'), -- i=717
      ("0101000101000000", '1'), -- i=718
      ("0100000101000000", '-'), -- i=719
      ("0000000111110100", '-'), -- i=720
      ("1000000101000111", '-'), -- i=721
      ("1001000101000111", '-'), -- i=722
      ("1010000101000111", '-'), -- i=723
      ("1011000101000111", '-'), -- i=724
      ("0101000101000000", '1'), -- i=725
      ("0100000101000000", '-'), -- i=726
      ("0000000110100101", '-'), -- i=727
      ("1000000101010000", '-'), -- i=728
      ("1001000101010000", '-'), -- i=729
      ("1010000101010000", '-'), -- i=730
      ("1011000101010000", '-'), -- i=731
      ("0101000101010000", '1'), -- i=732
      ("0100000101010000", '-'), -- i=733
      ("0000000110111111", '-'), -- i=734
      ("1000000101010001", '-'), -- i=735
      ("1001000101010001", '-'), -- i=736
      ("1010000101010001", '-'), -- i=737
      ("1011000101010001", '-'), -- i=738
      ("0101000101010000", '1'), -- i=739
      ("0100000101010000", '-'), -- i=740
      ("0000000111100010", '-'), -- i=741
      ("1000000101010010", '-'), -- i=742
      ("1001000101010010", '-'), -- i=743
      ("1010000101010010", '-'), -- i=744
      ("1011000101010010", '-'), -- i=745
      ("0101000101010000", '1'), -- i=746
      ("0100000101010000", '-'), -- i=747
      ("0000000100010010", '-'), -- i=748
      ("1000000101010011", '-'), -- i=749
      ("1001000101010011", '-'), -- i=750
      ("1010000101010011", '-'), -- i=751
      ("1011000101010011", '-'), -- i=752
      ("0101000101010000", '1'), -- i=753
      ("0100000101010000", '-'), -- i=754
      ("0000000111111001", '-'), -- i=755
      ("1000000101010100", '-'), -- i=756
      ("1001000101010100", '-'), -- i=757
      ("1010000101010100", '-'), -- i=758
      ("1011000101010100", '-'), -- i=759
      ("0101000101010000", '1'), -- i=760
      ("0100000101010000", '-'), -- i=761
      ("0000000101010111", '-'), -- i=762
      ("1000000101010101", '-'), -- i=763
      ("1001000101010101", '-'), -- i=764
      ("1010000101010101", '-'), -- i=765
      ("1011000101010101", '-'), -- i=766
      ("0101000101010000", '1'), -- i=767
      ("0100000101010000", '-'), -- i=768
      ("0000000111111000", '-'), -- i=769
      ("1000000101010110", '-'), -- i=770
      ("1001000101010110", '-'), -- i=771
      ("1010000101010110", '-'), -- i=772
      ("1011000101010110", '-'), -- i=773
      ("0101000101010000", '1'), -- i=774
      ("0100000101010000", '-'), -- i=775
      ("0000000111011010", '-'), -- i=776
      ("1000000101010111", '-'), -- i=777
      ("1001000101010111", '-'), -- i=778
      ("1010000101010111", '-'), -- i=779
      ("1011000101010111", '-'), -- i=780
      ("0101000101010000", '1'), -- i=781
      ("0100000101010000", '-'), -- i=782
      ("0000000100111101", '-'), -- i=783
      ("1000000101100000", '-'), -- i=784
      ("1001000101100000", '-'), -- i=785
      ("1010000101100000", '-'), -- i=786
      ("1011000101100000", '-'), -- i=787
      ("0101000101100000", '1'), -- i=788
      ("0100000101100000", '-'), -- i=789
      ("0000000101010010", '-'), -- i=790
      ("1000000101100001", '-'), -- i=791
      ("1001000101100001", '-'), -- i=792
      ("1010000101100001", '-'), -- i=793
      ("1011000101100001", '-'), -- i=794
      ("0101000101100000", '1'), -- i=795
      ("0100000101100000", '-'), -- i=796
      ("0000000111011001", '-'), -- i=797
      ("1000000101100010", '-'), -- i=798
      ("1001000101100010", '-'), -- i=799
      ("1010000101100010", '-'), -- i=800
      ("1011000101100010", '-'), -- i=801
      ("0101000101100000", '1'), -- i=802
      ("0100000101100000", '-'), -- i=803
      ("0000000111000111", '-'), -- i=804
      ("1000000101100011", '-'), -- i=805
      ("1001000101100011", '-'), -- i=806
      ("1010000101100011", '-'), -- i=807
      ("1011000101100011", '-'), -- i=808
      ("0101000101100000", '1'), -- i=809
      ("0100000101100000", '-'), -- i=810
      ("0000000101010001", '-'), -- i=811
      ("1000000101100100", '-'), -- i=812
      ("1001000101100100", '-'), -- i=813
      ("1010000101100100", '-'), -- i=814
      ("1011000101100100", '-'), -- i=815
      ("0101000101100000", '1'), -- i=816
      ("0100000101100000", '-'), -- i=817
      ("0000000101111111", '-'), -- i=818
      ("1000000101100101", '-'), -- i=819
      ("1001000101100101", '-'), -- i=820
      ("1010000101100101", '-'), -- i=821
      ("1011000101100101", '-'), -- i=822
      ("0101000101100000", '1'), -- i=823
      ("0100000101100000", '-'), -- i=824
      ("0000000111010001", '-'), -- i=825
      ("1000000101100110", '-'), -- i=826
      ("1001000101100110", '-'), -- i=827
      ("1010000101100110", '-'), -- i=828
      ("1011000101100110", '-'), -- i=829
      ("0101000101100000", '1'), -- i=830
      ("0100000101100000", '-'), -- i=831
      ("0000000101100010", '-'), -- i=832
      ("1000000101100111", '-'), -- i=833
      ("1001000101100111", '-'), -- i=834
      ("1010000101100111", '-'), -- i=835
      ("1011000101100111", '-'), -- i=836
      ("0101000101100000", '1'), -- i=837
      ("0100000101100000", '-'), -- i=838
      ("0000000100010110", '-'), -- i=839
      ("1000000101110000", '-'), -- i=840
      ("1001000101110000", '-'), -- i=841
      ("1010000101110000", '-'), -- i=842
      ("1011000101110000", '-'), -- i=843
      ("0101000101110000", '1'), -- i=844
      ("0100000101110000", '-'), -- i=845
      ("0000000110010101", '-'), -- i=846
      ("1000000101110001", '-'), -- i=847
      ("1001000101110001", '-'), -- i=848
      ("1010000101110001", '-'), -- i=849
      ("1011000101110001", '-'), -- i=850
      ("0101000101110000", '1'), -- i=851
      ("0100000101110000", '-'), -- i=852
      ("0000000100100101", '-'), -- i=853
      ("1000000101110010", '-'), -- i=854
      ("1001000101110010", '-'), -- i=855
      ("1010000101110010", '-'), -- i=856
      ("1011000101110010", '-'), -- i=857
      ("0101000101110000", '1'), -- i=858
      ("0100000101110000", '-'), -- i=859
      ("0000000100100001", '-'), -- i=860
      ("1000000101110011", '-'), -- i=861
      ("1001000101110011", '-'), -- i=862
      ("1010000101110011", '-'), -- i=863
      ("1011000101110011", '-'), -- i=864
      ("0101000101110000", '1'), -- i=865
      ("0100000101110000", '-'), -- i=866
      ("0000000110011000", '-'), -- i=867
      ("1000000101110100", '-'), -- i=868
      ("1001000101110100", '-'), -- i=869
      ("1010000101110100", '-'), -- i=870
      ("1011000101110100", '-'), -- i=871
      ("0101000101110000", '1'), -- i=872
      ("0100000101110000", '-'), -- i=873
      ("0000000110000000", '-'), -- i=874
      ("1000000101110101", '-'), -- i=875
      ("1001000101110101", '-'), -- i=876
      ("1010000101110101", '-'), -- i=877
      ("1011000101110101", '-'), -- i=878
      ("0101000101110000", '1'), -- i=879
      ("0100000101110000", '-'), -- i=880
      ("0000000100111110", '-'), -- i=881
      ("1000000101110110", '-'), -- i=882
      ("1001000101110110", '-'), -- i=883
      ("1010000101110110", '-'), -- i=884
      ("1011000101110110", '-'), -- i=885
      ("0101000101110000", '1'), -- i=886
      ("0100000101110000", '-'), -- i=887
      ("0000000100000010", '-'), -- i=888
      ("1000000101110111", '-'), -- i=889
      ("1001000101110111", '-'), -- i=890
      ("1010000101110111", '-'), -- i=891
      ("1011000101110111", '-'), -- i=892
      ("0101000101110000", '1'), -- i=893
      ("0100000101110000", '-'), -- i=894
      ("0000000111000010", '-'), -- i=895
      ("1000001000000000", '-'), -- i=896
      ("1001001000000000", '-'), -- i=897
      ("1010001000000000", '-'), -- i=898
      ("1011001000000000", '-'), -- i=899
      ("0101001000000000", '1'), -- i=900
      ("0100001000000000", '-'), -- i=901
      ("0000001000000010", '-'), -- i=902
      ("1000001000000001", '-'), -- i=903
      ("1001001000000001", '-'), -- i=904
      ("1010001000000001", '-'), -- i=905
      ("1011001000000001", '-'), -- i=906
      ("0101001000000000", '1'), -- i=907
      ("0100001000000000", '-'), -- i=908
      ("0000001011100001", '-'), -- i=909
      ("1000001000000010", '-'), -- i=910
      ("1001001000000010", '-'), -- i=911
      ("1010001000000010", '-'), -- i=912
      ("1011001000000010", '-'), -- i=913
      ("0101001000000000", '1'), -- i=914
      ("0100001000000000", '-'), -- i=915
      ("0000001011101000", '-'), -- i=916
      ("1000001000000011", '-'), -- i=917
      ("1001001000000011", '-'), -- i=918
      ("1010001000000011", '-'), -- i=919
      ("1011001000000011", '-'), -- i=920
      ("0101001000000000", '1'), -- i=921
      ("0100001000000000", '-'), -- i=922
      ("0000001001010010", '-'), -- i=923
      ("1000001000000100", '-'), -- i=924
      ("1001001000000100", '-'), -- i=925
      ("1010001000000100", '-'), -- i=926
      ("1011001000000100", '-'), -- i=927
      ("0101001000000000", '1'), -- i=928
      ("0100001000000000", '-'), -- i=929
      ("0000001001000111", '-'), -- i=930
      ("1000001000000101", '-'), -- i=931
      ("1001001000000101", '-'), -- i=932
      ("1010001000000101", '-'), -- i=933
      ("1011001000000101", '-'), -- i=934
      ("0101001000000000", '1'), -- i=935
      ("0100001000000000", '-'), -- i=936
      ("0000001011111101", '-'), -- i=937
      ("1000001000000110", '-'), -- i=938
      ("1001001000000110", '-'), -- i=939
      ("1010001000000110", '-'), -- i=940
      ("1011001000000110", '-'), -- i=941
      ("0101001000000000", '1'), -- i=942
      ("0100001000000000", '-'), -- i=943
      ("0000001001110001", '-'), -- i=944
      ("1000001000000111", '-'), -- i=945
      ("1001001000000111", '-'), -- i=946
      ("1010001000000111", '-'), -- i=947
      ("1011001000000111", '-'), -- i=948
      ("0101001000000000", '1'), -- i=949
      ("0100001000000000", '-'), -- i=950
      ("0000001010000111", '-'), -- i=951
      ("1000001000010000", '-'), -- i=952
      ("1001001000010000", '-'), -- i=953
      ("1010001000010000", '-'), -- i=954
      ("1011001000010000", '-'), -- i=955
      ("0101001000010000", '1'), -- i=956
      ("0100001000010000", '-'), -- i=957
      ("0000001011011111", '-'), -- i=958
      ("1000001000010001", '-'), -- i=959
      ("1001001000010001", '-'), -- i=960
      ("1010001000010001", '-'), -- i=961
      ("1011001000010001", '-'), -- i=962
      ("0101001000010000", '1'), -- i=963
      ("0100001000010000", '-'), -- i=964
      ("0000001011001010", '-'), -- i=965
      ("1000001000010010", '-'), -- i=966
      ("1001001000010010", '-'), -- i=967
      ("1010001000010010", '-'), -- i=968
      ("1011001000010010", '-'), -- i=969
      ("0101001000010000", '1'), -- i=970
      ("0100001000010000", '-'), -- i=971
      ("0000001000000111", '-'), -- i=972
      ("1000001000010011", '-'), -- i=973
      ("1001001000010011", '-'), -- i=974
      ("1010001000010011", '-'), -- i=975
      ("1011001000010011", '-'), -- i=976
      ("0101001000010000", '1'), -- i=977
      ("0100001000010000", '-'), -- i=978
      ("0000001011110000", '-'), -- i=979
      ("1000001000010100", '-'), -- i=980
      ("1001001000010100", '-'), -- i=981
      ("1010001000010100", '-'), -- i=982
      ("1011001000010100", '-'), -- i=983
      ("0101001000010000", '1'), -- i=984
      ("0100001000010000", '-'), -- i=985
      ("0000001010111110", '-'), -- i=986
      ("1000001000010101", '-'), -- i=987
      ("1001001000010101", '-'), -- i=988
      ("1010001000010101", '-'), -- i=989
      ("1011001000010101", '-'), -- i=990
      ("0101001000010000", '1'), -- i=991
      ("0100001000010000", '-'), -- i=992
      ("0000001000000111", '-'), -- i=993
      ("1000001000010110", '-'), -- i=994
      ("1001001000010110", '-'), -- i=995
      ("1010001000010110", '-'), -- i=996
      ("1011001000010110", '-'), -- i=997
      ("0101001000010000", '1'), -- i=998
      ("0100001000010000", '-'), -- i=999
      ("0000001010010110", '-'), -- i=1000
      ("1000001000010111", '-'), -- i=1001
      ("1001001000010111", '-'), -- i=1002
      ("1010001000010111", '-'), -- i=1003
      ("1011001000010111", '-'), -- i=1004
      ("0101001000010000", '1'), -- i=1005
      ("0100001000010000", '-'), -- i=1006
      ("0000001000111010", '-'), -- i=1007
      ("1000001000100000", '-'), -- i=1008
      ("1001001000100000", '-'), -- i=1009
      ("1010001000100000", '-'), -- i=1010
      ("1011001000100000", '-'), -- i=1011
      ("0101001000100000", '1'), -- i=1012
      ("0100001000100000", '-'), -- i=1013
      ("0000001010111000", '-'), -- i=1014
      ("1000001000100001", '-'), -- i=1015
      ("1001001000100001", '-'), -- i=1016
      ("1010001000100001", '-'), -- i=1017
      ("1011001000100001", '-'), -- i=1018
      ("0101001000100000", '1'), -- i=1019
      ("0100001000100000", '-'), -- i=1020
      ("0000001011010100", '-'), -- i=1021
      ("1000001000100010", '-'), -- i=1022
      ("1001001000100010", '-'), -- i=1023
      ("1010001000100010", '-'), -- i=1024
      ("1011001000100010", '-'), -- i=1025
      ("0101001000100000", '1'), -- i=1026
      ("0100001000100000", '-'), -- i=1027
      ("0000001001110011", '-'), -- i=1028
      ("1000001000100011", '-'), -- i=1029
      ("1001001000100011", '-'), -- i=1030
      ("1010001000100011", '-'), -- i=1031
      ("1011001000100011", '-'), -- i=1032
      ("0101001000100000", '1'), -- i=1033
      ("0100001000100000", '-'), -- i=1034
      ("0000001000111001", '-'), -- i=1035
      ("1000001000100100", '-'), -- i=1036
      ("1001001000100100", '-'), -- i=1037
      ("1010001000100100", '-'), -- i=1038
      ("1011001000100100", '-'), -- i=1039
      ("0101001000100000", '1'), -- i=1040
      ("0100001000100000", '-'), -- i=1041
      ("0000001000100011", '-'), -- i=1042
      ("1000001000100101", '-'), -- i=1043
      ("1001001000100101", '-'), -- i=1044
      ("1010001000100101", '-'), -- i=1045
      ("1011001000100101", '-'), -- i=1046
      ("0101001000100000", '1'), -- i=1047
      ("0100001000100000", '-'), -- i=1048
      ("0000001001110110", '-'), -- i=1049
      ("1000001000100110", '-'), -- i=1050
      ("1001001000100110", '-'), -- i=1051
      ("1010001000100110", '-'), -- i=1052
      ("1011001000100110", '-'), -- i=1053
      ("0101001000100000", '1'), -- i=1054
      ("0100001000100000", '-'), -- i=1055
      ("0000001011000101", '-'), -- i=1056
      ("1000001000100111", '-'), -- i=1057
      ("1001001000100111", '-'), -- i=1058
      ("1010001000100111", '-'), -- i=1059
      ("1011001000100111", '-'), -- i=1060
      ("0101001000100000", '1'), -- i=1061
      ("0100001000100000", '-'), -- i=1062
      ("0000001001111000", '-'), -- i=1063
      ("1000001000110000", '-'), -- i=1064
      ("1001001000110000", '-'), -- i=1065
      ("1010001000110000", '-'), -- i=1066
      ("1011001000110000", '-'), -- i=1067
      ("0101001000110000", '1'), -- i=1068
      ("0100001000110000", '-'), -- i=1069
      ("0000001001000100", '-'), -- i=1070
      ("1000001000110001", '-'), -- i=1071
      ("1001001000110001", '-'), -- i=1072
      ("1010001000110001", '-'), -- i=1073
      ("1011001000110001", '-'), -- i=1074
      ("0101001000110000", '1'), -- i=1075
      ("0100001000110000", '-'), -- i=1076
      ("0000001001110100", '-'), -- i=1077
      ("1000001000110010", '-'), -- i=1078
      ("1001001000110010", '-'), -- i=1079
      ("1010001000110010", '-'), -- i=1080
      ("1011001000110010", '-'), -- i=1081
      ("0101001000110000", '1'), -- i=1082
      ("0100001000110000", '-'), -- i=1083
      ("0000001011100110", '-'), -- i=1084
      ("1000001000110011", '-'), -- i=1085
      ("1001001000110011", '-'), -- i=1086
      ("1010001000110011", '-'), -- i=1087
      ("1011001000110011", '-'), -- i=1088
      ("0101001000110000", '1'), -- i=1089
      ("0100001000110000", '-'), -- i=1090
      ("0000001010011111", '-'), -- i=1091
      ("1000001000110100", '-'), -- i=1092
      ("1001001000110100", '-'), -- i=1093
      ("1010001000110100", '-'), -- i=1094
      ("1011001000110100", '-'), -- i=1095
      ("0101001000110000", '1'), -- i=1096
      ("0100001000110000", '-'), -- i=1097
      ("0000001001100111", '-'), -- i=1098
      ("1000001000110101", '-'), -- i=1099
      ("1001001000110101", '-'), -- i=1100
      ("1010001000110101", '-'), -- i=1101
      ("1011001000110101", '-'), -- i=1102
      ("0101001000110000", '1'), -- i=1103
      ("0100001000110000", '-'), -- i=1104
      ("0000001011011011", '-'), -- i=1105
      ("1000001000110110", '-'), -- i=1106
      ("1001001000110110", '-'), -- i=1107
      ("1010001000110110", '-'), -- i=1108
      ("1011001000110110", '-'), -- i=1109
      ("0101001000110000", '1'), -- i=1110
      ("0100001000110000", '-'), -- i=1111
      ("0000001011111110", '-'), -- i=1112
      ("1000001000110111", '-'), -- i=1113
      ("1001001000110111", '-'), -- i=1114
      ("1010001000110111", '-'), -- i=1115
      ("1011001000110111", '-'), -- i=1116
      ("0101001000110000", '1'), -- i=1117
      ("0100001000110000", '-'), -- i=1118
      ("0000001001101101", '-'), -- i=1119
      ("1000001001000000", '-'), -- i=1120
      ("1001001001000000", '-'), -- i=1121
      ("1010001001000000", '-'), -- i=1122
      ("1011001001000000", '-'), -- i=1123
      ("0101001001000000", '1'), -- i=1124
      ("0100001001000000", '-'), -- i=1125
      ("0000001001111001", '-'), -- i=1126
      ("1000001001000001", '-'), -- i=1127
      ("1001001001000001", '-'), -- i=1128
      ("1010001001000001", '-'), -- i=1129
      ("1011001001000001", '-'), -- i=1130
      ("0101001001000000", '1'), -- i=1131
      ("0100001001000000", '-'), -- i=1132
      ("0000001001000010", '-'), -- i=1133
      ("1000001001000010", '-'), -- i=1134
      ("1001001001000010", '-'), -- i=1135
      ("1010001001000010", '-'), -- i=1136
      ("1011001001000010", '-'), -- i=1137
      ("0101001001000000", '1'), -- i=1138
      ("0100001001000000", '-'), -- i=1139
      ("0000001001100111", '-'), -- i=1140
      ("1000001001000011", '-'), -- i=1141
      ("1001001001000011", '-'), -- i=1142
      ("1010001001000011", '-'), -- i=1143
      ("1011001001000011", '-'), -- i=1144
      ("0101001001000000", '1'), -- i=1145
      ("0100001001000000", '-'), -- i=1146
      ("0000001011010011", '-'), -- i=1147
      ("1000001001000100", '-'), -- i=1148
      ("1001001001000100", '-'), -- i=1149
      ("1010001001000100", '-'), -- i=1150
      ("1011001001000100", '-'), -- i=1151
      ("0101001001000000", '1'), -- i=1152
      ("0100001001000000", '-'), -- i=1153
      ("0000001001111010", '-'), -- i=1154
      ("1000001001000101", '-'), -- i=1155
      ("1001001001000101", '-'), -- i=1156
      ("1010001001000101", '-'), -- i=1157
      ("1011001001000101", '-'), -- i=1158
      ("0101001001000000", '1'), -- i=1159
      ("0100001001000000", '-'), -- i=1160
      ("0000001011110000", '-'), -- i=1161
      ("1000001001000110", '-'), -- i=1162
      ("1001001001000110", '-'), -- i=1163
      ("1010001001000110", '-'), -- i=1164
      ("1011001001000110", '-'), -- i=1165
      ("0101001001000000", '1'), -- i=1166
      ("0100001001000000", '-'), -- i=1167
      ("0000001000111001", '-'), -- i=1168
      ("1000001001000111", '-'), -- i=1169
      ("1001001001000111", '-'), -- i=1170
      ("1010001001000111", '-'), -- i=1171
      ("1011001001000111", '-'), -- i=1172
      ("0101001001000000", '1'), -- i=1173
      ("0100001001000000", '-'), -- i=1174
      ("0000001010010000", '-'), -- i=1175
      ("1000001001010000", '-'), -- i=1176
      ("1001001001010000", '-'), -- i=1177
      ("1010001001010000", '-'), -- i=1178
      ("1011001001010000", '-'), -- i=1179
      ("0101001001010000", '1'), -- i=1180
      ("0100001001010000", '-'), -- i=1181
      ("0000001011100000", '-'), -- i=1182
      ("1000001001010001", '-'), -- i=1183
      ("1001001001010001", '-'), -- i=1184
      ("1010001001010001", '-'), -- i=1185
      ("1011001001010001", '-'), -- i=1186
      ("0101001001010000", '1'), -- i=1187
      ("0100001001010000", '-'), -- i=1188
      ("0000001000000001", '-'), -- i=1189
      ("1000001001010010", '-'), -- i=1190
      ("1001001001010010", '-'), -- i=1191
      ("1010001001010010", '-'), -- i=1192
      ("1011001001010010", '-'), -- i=1193
      ("0101001001010000", '1'), -- i=1194
      ("0100001001010000", '-'), -- i=1195
      ("0000001010101010", '-'), -- i=1196
      ("1000001001010011", '-'), -- i=1197
      ("1001001001010011", '-'), -- i=1198
      ("1010001001010011", '-'), -- i=1199
      ("1011001001010011", '-'), -- i=1200
      ("0101001001010000", '1'), -- i=1201
      ("0100001001010000", '-'), -- i=1202
      ("0000001000011000", '-'), -- i=1203
      ("1000001001010100", '-'), -- i=1204
      ("1001001001010100", '-'), -- i=1205
      ("1010001001010100", '-'), -- i=1206
      ("1011001001010100", '-'), -- i=1207
      ("0101001001010000", '1'), -- i=1208
      ("0100001001010000", '-'), -- i=1209
      ("0000001011000100", '-'), -- i=1210
      ("1000001001010101", '-'), -- i=1211
      ("1001001001010101", '-'), -- i=1212
      ("1010001001010101", '-'), -- i=1213
      ("1011001001010101", '-'), -- i=1214
      ("0101001001010000", '1'), -- i=1215
      ("0100001001010000", '-'), -- i=1216
      ("0000001010111000", '-'), -- i=1217
      ("1000001001010110", '-'), -- i=1218
      ("1001001001010110", '-'), -- i=1219
      ("1010001001010110", '-'), -- i=1220
      ("1011001001010110", '-'), -- i=1221
      ("0101001001010000", '1'), -- i=1222
      ("0100001001010000", '-'), -- i=1223
      ("0000001011111010", '-'), -- i=1224
      ("1000001001010111", '-'), -- i=1225
      ("1001001001010111", '-'), -- i=1226
      ("1010001001010111", '-'), -- i=1227
      ("1011001001010111", '-'), -- i=1228
      ("0101001001010000", '1'), -- i=1229
      ("0100001001010000", '-'), -- i=1230
      ("0000001000000011", '-'), -- i=1231
      ("1000001001100000", '-'), -- i=1232
      ("1001001001100000", '-'), -- i=1233
      ("1010001001100000", '-'), -- i=1234
      ("1011001001100000", '-'), -- i=1235
      ("0101001001100000", '1'), -- i=1236
      ("0100001001100000", '-'), -- i=1237
      ("0000001010000011", '-'), -- i=1238
      ("1000001001100001", '-'), -- i=1239
      ("1001001001100001", '-'), -- i=1240
      ("1010001001100001", '-'), -- i=1241
      ("1011001001100001", '-'), -- i=1242
      ("0101001001100000", '1'), -- i=1243
      ("0100001001100000", '-'), -- i=1244
      ("0000001000101100", '-'), -- i=1245
      ("1000001001100010", '-'), -- i=1246
      ("1001001001100010", '-'), -- i=1247
      ("1010001001100010", '-'), -- i=1248
      ("1011001001100010", '-'), -- i=1249
      ("0101001001100000", '1'), -- i=1250
      ("0100001001100000", '-'), -- i=1251
      ("0000001010111101", '-'), -- i=1252
      ("1000001001100011", '-'), -- i=1253
      ("1001001001100011", '-'), -- i=1254
      ("1010001001100011", '-'), -- i=1255
      ("1011001001100011", '-'), -- i=1256
      ("0101001001100000", '1'), -- i=1257
      ("0100001001100000", '-'), -- i=1258
      ("0000001000100011", '-'), -- i=1259
      ("1000001001100100", '-'), -- i=1260
      ("1001001001100100", '-'), -- i=1261
      ("1010001001100100", '-'), -- i=1262
      ("1011001001100100", '-'), -- i=1263
      ("0101001001100000", '1'), -- i=1264
      ("0100001001100000", '-'), -- i=1265
      ("0000001000101001", '-'), -- i=1266
      ("1000001001100101", '-'), -- i=1267
      ("1001001001100101", '-'), -- i=1268
      ("1010001001100101", '-'), -- i=1269
      ("1011001001100101", '-'), -- i=1270
      ("0101001001100000", '1'), -- i=1271
      ("0100001001100000", '-'), -- i=1272
      ("0000001001100111", '-'), -- i=1273
      ("1000001001100110", '-'), -- i=1274
      ("1001001001100110", '-'), -- i=1275
      ("1010001001100110", '-'), -- i=1276
      ("1011001001100110", '-'), -- i=1277
      ("0101001001100000", '1'), -- i=1278
      ("0100001001100000", '-'), -- i=1279
      ("0000001010111001", '-'), -- i=1280
      ("1000001001100111", '-'), -- i=1281
      ("1001001001100111", '-'), -- i=1282
      ("1010001001100111", '-'), -- i=1283
      ("1011001001100111", '-'), -- i=1284
      ("0101001001100000", '1'), -- i=1285
      ("0100001001100000", '-'), -- i=1286
      ("0000001001111000", '-'), -- i=1287
      ("1000001001110000", '-'), -- i=1288
      ("1001001001110000", '-'), -- i=1289
      ("1010001001110000", '-'), -- i=1290
      ("1011001001110000", '-'), -- i=1291
      ("0101001001110000", '1'), -- i=1292
      ("0100001001110000", '-'), -- i=1293
      ("0000001000000010", '-'), -- i=1294
      ("1000001001110001", '-'), -- i=1295
      ("1001001001110001", '-'), -- i=1296
      ("1010001001110001", '-'), -- i=1297
      ("1011001001110001", '-'), -- i=1298
      ("0101001001110000", '1'), -- i=1299
      ("0100001001110000", '-'), -- i=1300
      ("0000001010100000", '-'), -- i=1301
      ("1000001001110010", '-'), -- i=1302
      ("1001001001110010", '-'), -- i=1303
      ("1010001001110010", '-'), -- i=1304
      ("1011001001110010", '-'), -- i=1305
      ("0101001001110000", '1'), -- i=1306
      ("0100001001110000", '-'), -- i=1307
      ("0000001010010000", '-'), -- i=1308
      ("1000001001110011", '-'), -- i=1309
      ("1001001001110011", '-'), -- i=1310
      ("1010001001110011", '-'), -- i=1311
      ("1011001001110011", '-'), -- i=1312
      ("0101001001110000", '1'), -- i=1313
      ("0100001001110000", '-'), -- i=1314
      ("0000001010010101", '-'), -- i=1315
      ("1000001001110100", '-'), -- i=1316
      ("1001001001110100", '-'), -- i=1317
      ("1010001001110100", '-'), -- i=1318
      ("1011001001110100", '-'), -- i=1319
      ("0101001001110000", '1'), -- i=1320
      ("0100001001110000", '-'), -- i=1321
      ("0000001001011110", '-'), -- i=1322
      ("1000001001110101", '-'), -- i=1323
      ("1001001001110101", '-'), -- i=1324
      ("1010001001110101", '-'), -- i=1325
      ("1011001001110101", '-'), -- i=1326
      ("0101001001110000", '1'), -- i=1327
      ("0100001001110000", '-'), -- i=1328
      ("0000001010101111", '-'), -- i=1329
      ("1000001001110110", '-'), -- i=1330
      ("1001001001110110", '-'), -- i=1331
      ("1010001001110110", '-'), -- i=1332
      ("1011001001110110", '-'), -- i=1333
      ("0101001001110000", '1'), -- i=1334
      ("0100001001110000", '-'), -- i=1335
      ("0000001011001110", '-'), -- i=1336
      ("1000001001110111", '-'), -- i=1337
      ("1001001001110111", '-'), -- i=1338
      ("1010001001110111", '-'), -- i=1339
      ("1011001001110111", '-'), -- i=1340
      ("0101001001110000", '1'), -- i=1341
      ("0100001001110000", '-'), -- i=1342
      ("0000001011001011", '-'), -- i=1343
      ("1000001100000000", '-'), -- i=1344
      ("1001001100000000", '-'), -- i=1345
      ("1010001100000000", '-'), -- i=1346
      ("1011001100000000", '-'), -- i=1347
      ("0101001100000000", '1'), -- i=1348
      ("0100001100000000", '-'), -- i=1349
      ("0000001110011101", '-'), -- i=1350
      ("1000001100000001", '-'), -- i=1351
      ("1001001100000001", '-'), -- i=1352
      ("1010001100000001", '-'), -- i=1353
      ("1011001100000001", '-'), -- i=1354
      ("0101001100000000", '1'), -- i=1355
      ("0100001100000000", '-'), -- i=1356
      ("0000001111111111", '-'), -- i=1357
      ("1000001100000010", '-'), -- i=1358
      ("1001001100000010", '-'), -- i=1359
      ("1010001100000010", '-'), -- i=1360
      ("1011001100000010", '-'), -- i=1361
      ("0101001100000000", '1'), -- i=1362
      ("0100001100000000", '-'), -- i=1363
      ("0000001101001001", '-'), -- i=1364
      ("1000001100000011", '-'), -- i=1365
      ("1001001100000011", '-'), -- i=1366
      ("1010001100000011", '-'), -- i=1367
      ("1011001100000011", '-'), -- i=1368
      ("0101001100000000", '1'), -- i=1369
      ("0100001100000000", '-'), -- i=1370
      ("0000001101001000", '-'), -- i=1371
      ("1000001100000100", '-'), -- i=1372
      ("1001001100000100", '-'), -- i=1373
      ("1010001100000100", '-'), -- i=1374
      ("1011001100000100", '-'), -- i=1375
      ("0101001100000000", '1'), -- i=1376
      ("0100001100000000", '-'), -- i=1377
      ("0000001101101111", '-'), -- i=1378
      ("1000001100000101", '-'), -- i=1379
      ("1001001100000101", '-'), -- i=1380
      ("1010001100000101", '-'), -- i=1381
      ("1011001100000101", '-'), -- i=1382
      ("0101001100000000", '1'), -- i=1383
      ("0100001100000000", '-'), -- i=1384
      ("0000001101000000", '-'), -- i=1385
      ("1000001100000110", '-'), -- i=1386
      ("1001001100000110", '-'), -- i=1387
      ("1010001100000110", '-'), -- i=1388
      ("1011001100000110", '-'), -- i=1389
      ("0101001100000000", '1'), -- i=1390
      ("0100001100000000", '-'), -- i=1391
      ("0000001111101100", '-'), -- i=1392
      ("1000001100000111", '-'), -- i=1393
      ("1001001100000111", '-'), -- i=1394
      ("1010001100000111", '-'), -- i=1395
      ("1011001100000111", '-'), -- i=1396
      ("0101001100000000", '1'), -- i=1397
      ("0100001100000000", '-'), -- i=1398
      ("0000001110101101", '-'), -- i=1399
      ("1000001100010000", '-'), -- i=1400
      ("1001001100010000", '-'), -- i=1401
      ("1010001100010000", '-'), -- i=1402
      ("1011001100010000", '-'), -- i=1403
      ("0101001100010000", '1'), -- i=1404
      ("0100001100010000", '-'), -- i=1405
      ("0000001101000010", '-'), -- i=1406
      ("1000001100010001", '-'), -- i=1407
      ("1001001100010001", '-'), -- i=1408
      ("1010001100010001", '-'), -- i=1409
      ("1011001100010001", '-'), -- i=1410
      ("0101001100010000", '1'), -- i=1411
      ("0100001100010000", '-'), -- i=1412
      ("0000001111010111", '-'), -- i=1413
      ("1000001100010010", '-'), -- i=1414
      ("1001001100010010", '-'), -- i=1415
      ("1010001100010010", '-'), -- i=1416
      ("1011001100010010", '-'), -- i=1417
      ("0101001100010000", '1'), -- i=1418
      ("0100001100010000", '-'), -- i=1419
      ("0000001110000000", '-'), -- i=1420
      ("1000001100010011", '-'), -- i=1421
      ("1001001100010011", '-'), -- i=1422
      ("1010001100010011", '-'), -- i=1423
      ("1011001100010011", '-'), -- i=1424
      ("0101001100010000", '1'), -- i=1425
      ("0100001100010000", '-'), -- i=1426
      ("0000001100001110", '-'), -- i=1427
      ("1000001100010100", '-'), -- i=1428
      ("1001001100010100", '-'), -- i=1429
      ("1010001100010100", '-'), -- i=1430
      ("1011001100010100", '-'), -- i=1431
      ("0101001100010000", '1'), -- i=1432
      ("0100001100010000", '-'), -- i=1433
      ("0000001110110000", '-'), -- i=1434
      ("1000001100010101", '-'), -- i=1435
      ("1001001100010101", '-'), -- i=1436
      ("1010001100010101", '-'), -- i=1437
      ("1011001100010101", '-'), -- i=1438
      ("0101001100010000", '1'), -- i=1439
      ("0100001100010000", '-'), -- i=1440
      ("0000001110011111", '-'), -- i=1441
      ("1000001100010110", '-'), -- i=1442
      ("1001001100010110", '-'), -- i=1443
      ("1010001100010110", '-'), -- i=1444
      ("1011001100010110", '-'), -- i=1445
      ("0101001100010000", '1'), -- i=1446
      ("0100001100010000", '-'), -- i=1447
      ("0000001101101111", '-'), -- i=1448
      ("1000001100010111", '-'), -- i=1449
      ("1001001100010111", '-'), -- i=1450
      ("1010001100010111", '-'), -- i=1451
      ("1011001100010111", '-'), -- i=1452
      ("0101001100010000", '1'), -- i=1453
      ("0100001100010000", '-'), -- i=1454
      ("0000001100100011", '-'), -- i=1455
      ("1000001100100000", '-'), -- i=1456
      ("1001001100100000", '-'), -- i=1457
      ("1010001100100000", '-'), -- i=1458
      ("1011001100100000", '-'), -- i=1459
      ("0101001100100000", '1'), -- i=1460
      ("0100001100100000", '-'), -- i=1461
      ("0000001111111110", '-'), -- i=1462
      ("1000001100100001", '-'), -- i=1463
      ("1001001100100001", '-'), -- i=1464
      ("1010001100100001", '-'), -- i=1465
      ("1011001100100001", '-'), -- i=1466
      ("0101001100100000", '1'), -- i=1467
      ("0100001100100000", '-'), -- i=1468
      ("0000001111000010", '-'), -- i=1469
      ("1000001100100010", '-'), -- i=1470
      ("1001001100100010", '-'), -- i=1471
      ("1010001100100010", '-'), -- i=1472
      ("1011001100100010", '-'), -- i=1473
      ("0101001100100000", '1'), -- i=1474
      ("0100001100100000", '-'), -- i=1475
      ("0000001110111001", '-'), -- i=1476
      ("1000001100100011", '-'), -- i=1477
      ("1001001100100011", '-'), -- i=1478
      ("1010001100100011", '-'), -- i=1479
      ("1011001100100011", '-'), -- i=1480
      ("0101001100100000", '1'), -- i=1481
      ("0100001100100000", '-'), -- i=1482
      ("0000001110011010", '-'), -- i=1483
      ("1000001100100100", '-'), -- i=1484
      ("1001001100100100", '-'), -- i=1485
      ("1010001100100100", '-'), -- i=1486
      ("1011001100100100", '-'), -- i=1487
      ("0101001100100000", '1'), -- i=1488
      ("0100001100100000", '-'), -- i=1489
      ("0000001110000111", '-'), -- i=1490
      ("1000001100100101", '-'), -- i=1491
      ("1001001100100101", '-'), -- i=1492
      ("1010001100100101", '-'), -- i=1493
      ("1011001100100101", '-'), -- i=1494
      ("0101001100100000", '1'), -- i=1495
      ("0100001100100000", '-'), -- i=1496
      ("0000001110101111", '-'), -- i=1497
      ("1000001100100110", '-'), -- i=1498
      ("1001001100100110", '-'), -- i=1499
      ("1010001100100110", '-'), -- i=1500
      ("1011001100100110", '-'), -- i=1501
      ("0101001100100000", '1'), -- i=1502
      ("0100001100100000", '-'), -- i=1503
      ("0000001111111100", '-'), -- i=1504
      ("1000001100100111", '-'), -- i=1505
      ("1001001100100111", '-'), -- i=1506
      ("1010001100100111", '-'), -- i=1507
      ("1011001100100111", '-'), -- i=1508
      ("0101001100100000", '1'), -- i=1509
      ("0100001100100000", '-'), -- i=1510
      ("0000001110100001", '-'), -- i=1511
      ("1000001100110000", '-'), -- i=1512
      ("1001001100110000", '-'), -- i=1513
      ("1010001100110000", '-'), -- i=1514
      ("1011001100110000", '-'), -- i=1515
      ("0101001100110000", '1'), -- i=1516
      ("0100001100110000", '-'), -- i=1517
      ("0000001101001111", '-'), -- i=1518
      ("1000001100110001", '-'), -- i=1519
      ("1001001100110001", '-'), -- i=1520
      ("1010001100110001", '-'), -- i=1521
      ("1011001100110001", '-'), -- i=1522
      ("0101001100110000", '1'), -- i=1523
      ("0100001100110000", '-'), -- i=1524
      ("0000001111110011", '-'), -- i=1525
      ("1000001100110010", '-'), -- i=1526
      ("1001001100110010", '-'), -- i=1527
      ("1010001100110010", '-'), -- i=1528
      ("1011001100110010", '-'), -- i=1529
      ("0101001100110000", '1'), -- i=1530
      ("0100001100110000", '-'), -- i=1531
      ("0000001111001110", '-'), -- i=1532
      ("1000001100110011", '-'), -- i=1533
      ("1001001100110011", '-'), -- i=1534
      ("1010001100110011", '-'), -- i=1535
      ("1011001100110011", '-'), -- i=1536
      ("0101001100110000", '1'), -- i=1537
      ("0100001100110000", '-'), -- i=1538
      ("0000001110100110", '-'), -- i=1539
      ("1000001100110100", '-'), -- i=1540
      ("1001001100110100", '-'), -- i=1541
      ("1010001100110100", '-'), -- i=1542
      ("1011001100110100", '-'), -- i=1543
      ("0101001100110000", '1'), -- i=1544
      ("0100001100110000", '-'), -- i=1545
      ("0000001111000011", '-'), -- i=1546
      ("1000001100110101", '-'), -- i=1547
      ("1001001100110101", '-'), -- i=1548
      ("1010001100110101", '-'), -- i=1549
      ("1011001100110101", '-'), -- i=1550
      ("0101001100110000", '1'), -- i=1551
      ("0100001100110000", '-'), -- i=1552
      ("0000001101110011", '-'), -- i=1553
      ("1000001100110110", '-'), -- i=1554
      ("1001001100110110", '-'), -- i=1555
      ("1010001100110110", '-'), -- i=1556
      ("1011001100110110", '-'), -- i=1557
      ("0101001100110000", '1'), -- i=1558
      ("0100001100110000", '-'), -- i=1559
      ("0000001100100101", '-'), -- i=1560
      ("1000001100110111", '-'), -- i=1561
      ("1001001100110111", '-'), -- i=1562
      ("1010001100110111", '-'), -- i=1563
      ("1011001100110111", '-'), -- i=1564
      ("0101001100110000", '1'), -- i=1565
      ("0100001100110000", '-'), -- i=1566
      ("0000001100000011", '-'), -- i=1567
      ("1000001101000000", '-'), -- i=1568
      ("1001001101000000", '-'), -- i=1569
      ("1010001101000000", '-'), -- i=1570
      ("1011001101000000", '-'), -- i=1571
      ("0101001101000000", '1'), -- i=1572
      ("0100001101000000", '-'), -- i=1573
      ("0000001100110110", '-'), -- i=1574
      ("1000001101000001", '-'), -- i=1575
      ("1001001101000001", '-'), -- i=1576
      ("1010001101000001", '-'), -- i=1577
      ("1011001101000001", '-'), -- i=1578
      ("0101001101000000", '1'), -- i=1579
      ("0100001101000000", '-'), -- i=1580
      ("0000001111110001", '-'), -- i=1581
      ("1000001101000010", '-'), -- i=1582
      ("1001001101000010", '-'), -- i=1583
      ("1010001101000010", '-'), -- i=1584
      ("1011001101000010", '-'), -- i=1585
      ("0101001101000000", '1'), -- i=1586
      ("0100001101000000", '-'), -- i=1587
      ("0000001100100101", '-'), -- i=1588
      ("1000001101000011", '-'), -- i=1589
      ("1001001101000011", '-'), -- i=1590
      ("1010001101000011", '-'), -- i=1591
      ("1011001101000011", '-'), -- i=1592
      ("0101001101000000", '1'), -- i=1593
      ("0100001101000000", '-'), -- i=1594
      ("0000001110010110", '-'), -- i=1595
      ("1000001101000100", '-'), -- i=1596
      ("1001001101000100", '-'), -- i=1597
      ("1010001101000100", '-'), -- i=1598
      ("1011001101000100", '-'), -- i=1599
      ("0101001101000000", '1'), -- i=1600
      ("0100001101000000", '-'), -- i=1601
      ("0000001101101001", '-'), -- i=1602
      ("1000001101000101", '-'), -- i=1603
      ("1001001101000101", '-'), -- i=1604
      ("1010001101000101", '-'), -- i=1605
      ("1011001101000101", '-'), -- i=1606
      ("0101001101000000", '1'), -- i=1607
      ("0100001101000000", '-'), -- i=1608
      ("0000001111111011", '-'), -- i=1609
      ("1000001101000110", '-'), -- i=1610
      ("1001001101000110", '-'), -- i=1611
      ("1010001101000110", '-'), -- i=1612
      ("1011001101000110", '-'), -- i=1613
      ("0101001101000000", '1'), -- i=1614
      ("0100001101000000", '-'), -- i=1615
      ("0000001100110001", '-'), -- i=1616
      ("1000001101000111", '-'), -- i=1617
      ("1001001101000111", '-'), -- i=1618
      ("1010001101000111", '-'), -- i=1619
      ("1011001101000111", '-'), -- i=1620
      ("0101001101000000", '1'), -- i=1621
      ("0100001101000000", '-'), -- i=1622
      ("0000001111000101", '-'), -- i=1623
      ("1000001101010000", '-'), -- i=1624
      ("1001001101010000", '-'), -- i=1625
      ("1010001101010000", '-'), -- i=1626
      ("1011001101010000", '-'), -- i=1627
      ("0101001101010000", '1'), -- i=1628
      ("0100001101010000", '-'), -- i=1629
      ("0000001100010011", '-'), -- i=1630
      ("1000001101010001", '-'), -- i=1631
      ("1001001101010001", '-'), -- i=1632
      ("1010001101010001", '-'), -- i=1633
      ("1011001101010001", '-'), -- i=1634
      ("0101001101010000", '1'), -- i=1635
      ("0100001101010000", '-'), -- i=1636
      ("0000001101110001", '-'), -- i=1637
      ("1000001101010010", '-'), -- i=1638
      ("1001001101010010", '-'), -- i=1639
      ("1010001101010010", '-'), -- i=1640
      ("1011001101010010", '-'), -- i=1641
      ("0101001101010000", '1'), -- i=1642
      ("0100001101010000", '-'), -- i=1643
      ("0000001111000100", '-'), -- i=1644
      ("1000001101010011", '-'), -- i=1645
      ("1001001101010011", '-'), -- i=1646
      ("1010001101010011", '-'), -- i=1647
      ("1011001101010011", '-'), -- i=1648
      ("0101001101010000", '1'), -- i=1649
      ("0100001101010000", '-'), -- i=1650
      ("0000001100101001", '-'), -- i=1651
      ("1000001101010100", '-'), -- i=1652
      ("1001001101010100", '-'), -- i=1653
      ("1010001101010100", '-'), -- i=1654
      ("1011001101010100", '-'), -- i=1655
      ("0101001101010000", '1'), -- i=1656
      ("0100001101010000", '-'), -- i=1657
      ("0000001100110100", '-'), -- i=1658
      ("1000001101010101", '-'), -- i=1659
      ("1001001101010101", '-'), -- i=1660
      ("1010001101010101", '-'), -- i=1661
      ("1011001101010101", '-'), -- i=1662
      ("0101001101010000", '1'), -- i=1663
      ("0100001101010000", '-'), -- i=1664
      ("0000001101111110", '-'), -- i=1665
      ("1000001101010110", '-'), -- i=1666
      ("1001001101010110", '-'), -- i=1667
      ("1010001101010110", '-'), -- i=1668
      ("1011001101010110", '-'), -- i=1669
      ("0101001101010000", '1'), -- i=1670
      ("0100001101010000", '-'), -- i=1671
      ("0000001100100101", '-'), -- i=1672
      ("1000001101010111", '-'), -- i=1673
      ("1001001101010111", '-'), -- i=1674
      ("1010001101010111", '-'), -- i=1675
      ("1011001101010111", '-'), -- i=1676
      ("0101001101010000", '1'), -- i=1677
      ("0100001101010000", '-'), -- i=1678
      ("0000001100100000", '-'), -- i=1679
      ("1000001101100000", '-'), -- i=1680
      ("1001001101100000", '-'), -- i=1681
      ("1010001101100000", '-'), -- i=1682
      ("1011001101100000", '-'), -- i=1683
      ("0101001101100000", '1'), -- i=1684
      ("0100001101100000", '-'), -- i=1685
      ("0000001110100001", '-'), -- i=1686
      ("1000001101100001", '-'), -- i=1687
      ("1001001101100001", '-'), -- i=1688
      ("1010001101100001", '-'), -- i=1689
      ("1011001101100001", '-'), -- i=1690
      ("0101001101100000", '1'), -- i=1691
      ("0100001101100000", '-'), -- i=1692
      ("0000001110001111", '-'), -- i=1693
      ("1000001101100010", '-'), -- i=1694
      ("1001001101100010", '-'), -- i=1695
      ("1010001101100010", '-'), -- i=1696
      ("1011001101100010", '-'), -- i=1697
      ("0101001101100000", '1'), -- i=1698
      ("0100001101100000", '-'), -- i=1699
      ("0000001111000010", '-'), -- i=1700
      ("1000001101100011", '-'), -- i=1701
      ("1001001101100011", '-'), -- i=1702
      ("1010001101100011", '-'), -- i=1703
      ("1011001101100011", '-'), -- i=1704
      ("0101001101100000", '1'), -- i=1705
      ("0100001101100000", '-'), -- i=1706
      ("0000001111111110", '-'), -- i=1707
      ("1000001101100100", '-'), -- i=1708
      ("1001001101100100", '-'), -- i=1709
      ("1010001101100100", '-'), -- i=1710
      ("1011001101100100", '-'), -- i=1711
      ("0101001101100000", '1'), -- i=1712
      ("0100001101100000", '-'), -- i=1713
      ("0000001100110001", '-'), -- i=1714
      ("1000001101100101", '-'), -- i=1715
      ("1001001101100101", '-'), -- i=1716
      ("1010001101100101", '-'), -- i=1717
      ("1011001101100101", '-'), -- i=1718
      ("0101001101100000", '1'), -- i=1719
      ("0100001101100000", '-'), -- i=1720
      ("0000001100001011", '-'), -- i=1721
      ("1000001101100110", '-'), -- i=1722
      ("1001001101100110", '-'), -- i=1723
      ("1010001101100110", '-'), -- i=1724
      ("1011001101100110", '-'), -- i=1725
      ("0101001101100000", '1'), -- i=1726
      ("0100001101100000", '-'), -- i=1727
      ("0000001110110010", '-'), -- i=1728
      ("1000001101100111", '-'), -- i=1729
      ("1001001101100111", '-'), -- i=1730
      ("1010001101100111", '-'), -- i=1731
      ("1011001101100111", '-'), -- i=1732
      ("0101001101100000", '1'), -- i=1733
      ("0100001101100000", '-'), -- i=1734
      ("0000001111110111", '-'), -- i=1735
      ("1000001101110000", '-'), -- i=1736
      ("1001001101110000", '-'), -- i=1737
      ("1010001101110000", '-'), -- i=1738
      ("1011001101110000", '-'), -- i=1739
      ("0101001101110000", '1'), -- i=1740
      ("0100001101110000", '-'), -- i=1741
      ("0000001110011011", '-'), -- i=1742
      ("1000001101110001", '-'), -- i=1743
      ("1001001101110001", '-'), -- i=1744
      ("1010001101110001", '-'), -- i=1745
      ("1011001101110001", '-'), -- i=1746
      ("0101001101110000", '1'), -- i=1747
      ("0100001101110000", '-'), -- i=1748
      ("0000001111010111", '-'), -- i=1749
      ("1000001101110010", '-'), -- i=1750
      ("1001001101110010", '-'), -- i=1751
      ("1010001101110010", '-'), -- i=1752
      ("1011001101110010", '-'), -- i=1753
      ("0101001101110000", '1'), -- i=1754
      ("0100001101110000", '-'), -- i=1755
      ("0000001110010001", '-'), -- i=1756
      ("1000001101110011", '-'), -- i=1757
      ("1001001101110011", '-'), -- i=1758
      ("1010001101110011", '-'), -- i=1759
      ("1011001101110011", '-'), -- i=1760
      ("0101001101110000", '1'), -- i=1761
      ("0100001101110000", '-'), -- i=1762
      ("0000001111111001", '-'), -- i=1763
      ("1000001101110100", '-'), -- i=1764
      ("1001001101110100", '-'), -- i=1765
      ("1010001101110100", '-'), -- i=1766
      ("1011001101110100", '-'), -- i=1767
      ("0101001101110000", '1'), -- i=1768
      ("0100001101110000", '-'), -- i=1769
      ("0000001100100100", '-'), -- i=1770
      ("1000001101110101", '-'), -- i=1771
      ("1001001101110101", '-'), -- i=1772
      ("1010001101110101", '-'), -- i=1773
      ("1011001101110101", '-'), -- i=1774
      ("0101001101110000", '1'), -- i=1775
      ("0100001101110000", '-'), -- i=1776
      ("0000001101100000", '-'), -- i=1777
      ("1000001101110110", '-'), -- i=1778
      ("1001001101110110", '-'), -- i=1779
      ("1010001101110110", '-'), -- i=1780
      ("1011001101110110", '-'), -- i=1781
      ("0101001101110000", '1'), -- i=1782
      ("0100001101110000", '-'), -- i=1783
      ("0000001110100111", '-'), -- i=1784
      ("1000001101110111", '-'), -- i=1785
      ("1001001101110111", '-'), -- i=1786
      ("1010001101110111", '-'), -- i=1787
      ("1011001101110111", '-'), -- i=1788
      ("0101001101110000", '1'), -- i=1789
      ("0100001101110000", '-'), -- i=1790
      ("0000001110111101", '-'), -- i=1791
      ("1000010000000000", '-'), -- i=1792
      ("1001010000000000", '-'), -- i=1793
      ("1010010000000000", '-'), -- i=1794
      ("1011010000000000", '-'), -- i=1795
      ("0101010000000000", '1'), -- i=1796
      ("0100010000000000", '-'), -- i=1797
      ("0000010011100110", '-'), -- i=1798
      ("1000010000000001", '-'), -- i=1799
      ("1001010000000001", '-'), -- i=1800
      ("1010010000000001", '-'), -- i=1801
      ("1011010000000001", '-'), -- i=1802
      ("0101010000000000", '1'), -- i=1803
      ("0100010000000000", '-'), -- i=1804
      ("0000010011100010", '-'), -- i=1805
      ("1000010000000010", '-'), -- i=1806
      ("1001010000000010", '-'), -- i=1807
      ("1010010000000010", '-'), -- i=1808
      ("1011010000000010", '-'), -- i=1809
      ("0101010000000000", '1'), -- i=1810
      ("0100010000000000", '-'), -- i=1811
      ("0000010000100110", '-'), -- i=1812
      ("1000010000000011", '-'), -- i=1813
      ("1001010000000011", '-'), -- i=1814
      ("1010010000000011", '-'), -- i=1815
      ("1011010000000011", '-'), -- i=1816
      ("0101010000000000", '1'), -- i=1817
      ("0100010000000000", '-'), -- i=1818
      ("0000010011000100", '-'), -- i=1819
      ("1000010000000100", '-'), -- i=1820
      ("1001010000000100", '-'), -- i=1821
      ("1010010000000100", '-'), -- i=1822
      ("1011010000000100", '-'), -- i=1823
      ("0101010000000000", '1'), -- i=1824
      ("0100010000000000", '-'), -- i=1825
      ("0000010010110110", '-'), -- i=1826
      ("1000010000000101", '-'), -- i=1827
      ("1001010000000101", '-'), -- i=1828
      ("1010010000000101", '-'), -- i=1829
      ("1011010000000101", '-'), -- i=1830
      ("0101010000000000", '1'), -- i=1831
      ("0100010000000000", '-'), -- i=1832
      ("0000010011000101", '-'), -- i=1833
      ("1000010000000110", '-'), -- i=1834
      ("1001010000000110", '-'), -- i=1835
      ("1010010000000110", '-'), -- i=1836
      ("1011010000000110", '-'), -- i=1837
      ("0101010000000000", '1'), -- i=1838
      ("0100010000000000", '-'), -- i=1839
      ("0000010000001001", '-'), -- i=1840
      ("1000010000000111", '-'), -- i=1841
      ("1001010000000111", '-'), -- i=1842
      ("1010010000000111", '-'), -- i=1843
      ("1011010000000111", '-'), -- i=1844
      ("0101010000000000", '1'), -- i=1845
      ("0100010000000000", '-'), -- i=1846
      ("0000010011000110", '-'), -- i=1847
      ("1000010000010000", '-'), -- i=1848
      ("1001010000010000", '-'), -- i=1849
      ("1010010000010000", '-'), -- i=1850
      ("1011010000010000", '-'), -- i=1851
      ("0101010000010000", '1'), -- i=1852
      ("0100010000010000", '-'), -- i=1853
      ("0000010001000111", '-'), -- i=1854
      ("1000010000010001", '-'), -- i=1855
      ("1001010000010001", '-'), -- i=1856
      ("1010010000010001", '-'), -- i=1857
      ("1011010000010001", '-'), -- i=1858
      ("0101010000010000", '1'), -- i=1859
      ("0100010000010000", '-'), -- i=1860
      ("0000010001110111", '-'), -- i=1861
      ("1000010000010010", '-'), -- i=1862
      ("1001010000010010", '-'), -- i=1863
      ("1010010000010010", '-'), -- i=1864
      ("1011010000010010", '-'), -- i=1865
      ("0101010000010000", '1'), -- i=1866
      ("0100010000010000", '-'), -- i=1867
      ("0000010000001000", '-'), -- i=1868
      ("1000010000010011", '-'), -- i=1869
      ("1001010000010011", '-'), -- i=1870
      ("1010010000010011", '-'), -- i=1871
      ("1011010000010011", '-'), -- i=1872
      ("0101010000010000", '1'), -- i=1873
      ("0100010000010000", '-'), -- i=1874
      ("0000010000001101", '-'), -- i=1875
      ("1000010000010100", '-'), -- i=1876
      ("1001010000010100", '-'), -- i=1877
      ("1010010000010100", '-'), -- i=1878
      ("1011010000010100", '-'), -- i=1879
      ("0101010000010000", '1'), -- i=1880
      ("0100010000010000", '-'), -- i=1881
      ("0000010010001100", '-'), -- i=1882
      ("1000010000010101", '-'), -- i=1883
      ("1001010000010101", '-'), -- i=1884
      ("1010010000010101", '-'), -- i=1885
      ("1011010000010101", '-'), -- i=1886
      ("0101010000010000", '1'), -- i=1887
      ("0100010000010000", '-'), -- i=1888
      ("0000010011111111", '-'), -- i=1889
      ("1000010000010110", '-'), -- i=1890
      ("1001010000010110", '-'), -- i=1891
      ("1010010000010110", '-'), -- i=1892
      ("1011010000010110", '-'), -- i=1893
      ("0101010000010000", '1'), -- i=1894
      ("0100010000010000", '-'), -- i=1895
      ("0000010011110011", '-'), -- i=1896
      ("1000010000010111", '-'), -- i=1897
      ("1001010000010111", '-'), -- i=1898
      ("1010010000010111", '-'), -- i=1899
      ("1011010000010111", '-'), -- i=1900
      ("0101010000010000", '1'), -- i=1901
      ("0100010000010000", '-'), -- i=1902
      ("0000010010010011", '-'), -- i=1903
      ("1000010000100000", '-'), -- i=1904
      ("1001010000100000", '-'), -- i=1905
      ("1010010000100000", '-'), -- i=1906
      ("1011010000100000", '-'), -- i=1907
      ("0101010000100000", '1'), -- i=1908
      ("0100010000100000", '-'), -- i=1909
      ("0000010011111100", '-'), -- i=1910
      ("1000010000100001", '-'), -- i=1911
      ("1001010000100001", '-'), -- i=1912
      ("1010010000100001", '-'), -- i=1913
      ("1011010000100001", '-'), -- i=1914
      ("0101010000100000", '1'), -- i=1915
      ("0100010000100000", '-'), -- i=1916
      ("0000010001101000", '-'), -- i=1917
      ("1000010000100010", '-'), -- i=1918
      ("1001010000100010", '-'), -- i=1919
      ("1010010000100010", '-'), -- i=1920
      ("1011010000100010", '-'), -- i=1921
      ("0101010000100000", '1'), -- i=1922
      ("0100010000100000", '-'), -- i=1923
      ("0000010010101010", '-'), -- i=1924
      ("1000010000100011", '-'), -- i=1925
      ("1001010000100011", '-'), -- i=1926
      ("1010010000100011", '-'), -- i=1927
      ("1011010000100011", '-'), -- i=1928
      ("0101010000100000", '1'), -- i=1929
      ("0100010000100000", '-'), -- i=1930
      ("0000010000101111", '-'), -- i=1931
      ("1000010000100100", '-'), -- i=1932
      ("1001010000100100", '-'), -- i=1933
      ("1010010000100100", '-'), -- i=1934
      ("1011010000100100", '-'), -- i=1935
      ("0101010000100000", '1'), -- i=1936
      ("0100010000100000", '-'), -- i=1937
      ("0000010011000100", '-'), -- i=1938
      ("1000010000100101", '-'), -- i=1939
      ("1001010000100101", '-'), -- i=1940
      ("1010010000100101", '-'), -- i=1941
      ("1011010000100101", '-'), -- i=1942
      ("0101010000100000", '1'), -- i=1943
      ("0100010000100000", '-'), -- i=1944
      ("0000010010111101", '-'), -- i=1945
      ("1000010000100110", '-'), -- i=1946
      ("1001010000100110", '-'), -- i=1947
      ("1010010000100110", '-'), -- i=1948
      ("1011010000100110", '-'), -- i=1949
      ("0101010000100000", '1'), -- i=1950
      ("0100010000100000", '-'), -- i=1951
      ("0000010011011100", '-'), -- i=1952
      ("1000010000100111", '-'), -- i=1953
      ("1001010000100111", '-'), -- i=1954
      ("1010010000100111", '-'), -- i=1955
      ("1011010000100111", '-'), -- i=1956
      ("0101010000100000", '1'), -- i=1957
      ("0100010000100000", '-'), -- i=1958
      ("0000010000100100", '-'), -- i=1959
      ("1000010000110000", '-'), -- i=1960
      ("1001010000110000", '-'), -- i=1961
      ("1010010000110000", '-'), -- i=1962
      ("1011010000110000", '-'), -- i=1963
      ("0101010000110000", '1'), -- i=1964
      ("0100010000110000", '-'), -- i=1965
      ("0000010011000100", '-'), -- i=1966
      ("1000010000110001", '-'), -- i=1967
      ("1001010000110001", '-'), -- i=1968
      ("1010010000110001", '-'), -- i=1969
      ("1011010000110001", '-'), -- i=1970
      ("0101010000110000", '1'), -- i=1971
      ("0100010000110000", '-'), -- i=1972
      ("0000010010101101", '-'), -- i=1973
      ("1000010000110010", '-'), -- i=1974
      ("1001010000110010", '-'), -- i=1975
      ("1010010000110010", '-'), -- i=1976
      ("1011010000110010", '-'), -- i=1977
      ("0101010000110000", '1'), -- i=1978
      ("0100010000110000", '-'), -- i=1979
      ("0000010011000001", '-'), -- i=1980
      ("1000010000110011", '-'), -- i=1981
      ("1001010000110011", '-'), -- i=1982
      ("1010010000110011", '-'), -- i=1983
      ("1011010000110011", '-'), -- i=1984
      ("0101010000110000", '1'), -- i=1985
      ("0100010000110000", '-'), -- i=1986
      ("0000010001100101", '-'), -- i=1987
      ("1000010000110100", '-'), -- i=1988
      ("1001010000110100", '-'), -- i=1989
      ("1010010000110100", '-'), -- i=1990
      ("1011010000110100", '-'), -- i=1991
      ("0101010000110000", '1'), -- i=1992
      ("0100010000110000", '-'), -- i=1993
      ("0000010010000010", '-'), -- i=1994
      ("1000010000110101", '-'), -- i=1995
      ("1001010000110101", '-'), -- i=1996
      ("1010010000110101", '-'), -- i=1997
      ("1011010000110101", '-'), -- i=1998
      ("0101010000110000", '1'), -- i=1999
      ("0100010000110000", '-'), -- i=2000
      ("0000010000001110", '-'), -- i=2001
      ("1000010000110110", '-'), -- i=2002
      ("1001010000110110", '-'), -- i=2003
      ("1010010000110110", '-'), -- i=2004
      ("1011010000110110", '-'), -- i=2005
      ("0101010000110000", '1'), -- i=2006
      ("0100010000110000", '-'), -- i=2007
      ("0000010011101001", '-'), -- i=2008
      ("1000010000110111", '-'), -- i=2009
      ("1001010000110111", '-'), -- i=2010
      ("1010010000110111", '-'), -- i=2011
      ("1011010000110111", '-'), -- i=2012
      ("0101010000110000", '1'), -- i=2013
      ("0100010000110000", '-'), -- i=2014
      ("0000010001011100", '-'), -- i=2015
      ("1000010001000000", '-'), -- i=2016
      ("1001010001000000", '-'), -- i=2017
      ("1010010001000000", '-'), -- i=2018
      ("1011010001000000", '-'), -- i=2019
      ("0101010001000000", '1'), -- i=2020
      ("0100010001000000", '-'), -- i=2021
      ("0000010000110101", '-'), -- i=2022
      ("1000010001000001", '-'), -- i=2023
      ("1001010001000001", '-'), -- i=2024
      ("1010010001000001", '-'), -- i=2025
      ("1011010001000001", '-'), -- i=2026
      ("0101010001000000", '1'), -- i=2027
      ("0100010001000000", '-'), -- i=2028
      ("0000010001110010", '-'), -- i=2029
      ("1000010001000010", '-'), -- i=2030
      ("1001010001000010", '-'), -- i=2031
      ("1010010001000010", '-'), -- i=2032
      ("1011010001000010", '-'), -- i=2033
      ("0101010001000000", '1'), -- i=2034
      ("0100010001000000", '-'), -- i=2035
      ("0000010001100000", '-'), -- i=2036
      ("1000010001000011", '-'), -- i=2037
      ("1001010001000011", '-'), -- i=2038
      ("1010010001000011", '-'), -- i=2039
      ("1011010001000011", '-'), -- i=2040
      ("0101010001000000", '1'), -- i=2041
      ("0100010001000000", '-'), -- i=2042
      ("0000010011000011", '-'), -- i=2043
      ("1000010001000100", '-'), -- i=2044
      ("1001010001000100", '-'), -- i=2045
      ("1010010001000100", '-'), -- i=2046
      ("1011010001000100", '-'), -- i=2047
      ("0101010001000000", '1'), -- i=2048
      ("0100010001000000", '-'), -- i=2049
      ("0000010010000001", '-'), -- i=2050
      ("1000010001000101", '-'), -- i=2051
      ("1001010001000101", '-'), -- i=2052
      ("1010010001000101", '-'), -- i=2053
      ("1011010001000101", '-'), -- i=2054
      ("0101010001000000", '1'), -- i=2055
      ("0100010001000000", '-'), -- i=2056
      ("0000010010111100", '-'), -- i=2057
      ("1000010001000110", '-'), -- i=2058
      ("1001010001000110", '-'), -- i=2059
      ("1010010001000110", '-'), -- i=2060
      ("1011010001000110", '-'), -- i=2061
      ("0101010001000000", '1'), -- i=2062
      ("0100010001000000", '-'), -- i=2063
      ("0000010001100011", '-'), -- i=2064
      ("1000010001000111", '-'), -- i=2065
      ("1001010001000111", '-'), -- i=2066
      ("1010010001000111", '-'), -- i=2067
      ("1011010001000111", '-'), -- i=2068
      ("0101010001000000", '1'), -- i=2069
      ("0100010001000000", '-'), -- i=2070
      ("0000010011110001", '-'), -- i=2071
      ("1000010001010000", '-'), -- i=2072
      ("1001010001010000", '-'), -- i=2073
      ("1010010001010000", '-'), -- i=2074
      ("1011010001010000", '-'), -- i=2075
      ("0101010001010000", '1'), -- i=2076
      ("0100010001010000", '-'), -- i=2077
      ("0000010001010001", '-'), -- i=2078
      ("1000010001010001", '-'), -- i=2079
      ("1001010001010001", '-'), -- i=2080
      ("1010010001010001", '-'), -- i=2081
      ("1011010001010001", '-'), -- i=2082
      ("0101010001010000", '1'), -- i=2083
      ("0100010001010000", '-'), -- i=2084
      ("0000010000001000", '-'), -- i=2085
      ("1000010001010010", '-'), -- i=2086
      ("1001010001010010", '-'), -- i=2087
      ("1010010001010010", '-'), -- i=2088
      ("1011010001010010", '-'), -- i=2089
      ("0101010001010000", '1'), -- i=2090
      ("0100010001010000", '-'), -- i=2091
      ("0000010000001101", '-'), -- i=2092
      ("1000010001010011", '-'), -- i=2093
      ("1001010001010011", '-'), -- i=2094
      ("1010010001010011", '-'), -- i=2095
      ("1011010001010011", '-'), -- i=2096
      ("0101010001010000", '1'), -- i=2097
      ("0100010001010000", '-'), -- i=2098
      ("0000010010000011", '-'), -- i=2099
      ("1000010001010100", '-'), -- i=2100
      ("1001010001010100", '-'), -- i=2101
      ("1010010001010100", '-'), -- i=2102
      ("1011010001010100", '-'), -- i=2103
      ("0101010001010000", '1'), -- i=2104
      ("0100010001010000", '-'), -- i=2105
      ("0000010011011101", '-'), -- i=2106
      ("1000010001010101", '-'), -- i=2107
      ("1001010001010101", '-'), -- i=2108
      ("1010010001010101", '-'), -- i=2109
      ("1011010001010101", '-'), -- i=2110
      ("0101010001010000", '1'), -- i=2111
      ("0100010001010000", '-'), -- i=2112
      ("0000010010101011", '-'), -- i=2113
      ("1000010001010110", '-'), -- i=2114
      ("1001010001010110", '-'), -- i=2115
      ("1010010001010110", '-'), -- i=2116
      ("1011010001010110", '-'), -- i=2117
      ("0101010001010000", '1'), -- i=2118
      ("0100010001010000", '-'), -- i=2119
      ("0000010001111111", '-'), -- i=2120
      ("1000010001010111", '-'), -- i=2121
      ("1001010001010111", '-'), -- i=2122
      ("1010010001010111", '-'), -- i=2123
      ("1011010001010111", '-'), -- i=2124
      ("0101010001010000", '1'), -- i=2125
      ("0100010001010000", '-'), -- i=2126
      ("0000010010000111", '-'), -- i=2127
      ("1000010001100000", '-'), -- i=2128
      ("1001010001100000", '-'), -- i=2129
      ("1010010001100000", '-'), -- i=2130
      ("1011010001100000", '-'), -- i=2131
      ("0101010001100000", '1'), -- i=2132
      ("0100010001100000", '-'), -- i=2133
      ("0000010011011011", '-'), -- i=2134
      ("1000010001100001", '-'), -- i=2135
      ("1001010001100001", '-'), -- i=2136
      ("1010010001100001", '-'), -- i=2137
      ("1011010001100001", '-'), -- i=2138
      ("0101010001100000", '1'), -- i=2139
      ("0100010001100000", '-'), -- i=2140
      ("0000010011111111", '-'), -- i=2141
      ("1000010001100010", '-'), -- i=2142
      ("1001010001100010", '-'), -- i=2143
      ("1010010001100010", '-'), -- i=2144
      ("1011010001100010", '-'), -- i=2145
      ("0101010001100000", '1'), -- i=2146
      ("0100010001100000", '-'), -- i=2147
      ("0000010000100111", '-'), -- i=2148
      ("1000010001100011", '-'), -- i=2149
      ("1001010001100011", '-'), -- i=2150
      ("1010010001100011", '-'), -- i=2151
      ("1011010001100011", '-'), -- i=2152
      ("0101010001100000", '1'), -- i=2153
      ("0100010001100000", '-'), -- i=2154
      ("0000010001101110", '-'), -- i=2155
      ("1000010001100100", '-'), -- i=2156
      ("1001010001100100", '-'), -- i=2157
      ("1010010001100100", '-'), -- i=2158
      ("1011010001100100", '-'), -- i=2159
      ("0101010001100000", '1'), -- i=2160
      ("0100010001100000", '-'), -- i=2161
      ("0000010001111011", '-'), -- i=2162
      ("1000010001100101", '-'), -- i=2163
      ("1001010001100101", '-'), -- i=2164
      ("1010010001100101", '-'), -- i=2165
      ("1011010001100101", '-'), -- i=2166
      ("0101010001100000", '1'), -- i=2167
      ("0100010001100000", '-'), -- i=2168
      ("0000010010001110", '-'), -- i=2169
      ("1000010001100110", '-'), -- i=2170
      ("1001010001100110", '-'), -- i=2171
      ("1010010001100110", '-'), -- i=2172
      ("1011010001100110", '-'), -- i=2173
      ("0101010001100000", '1'), -- i=2174
      ("0100010001100000", '-'), -- i=2175
      ("0000010000001101", '-'), -- i=2176
      ("1000010001100111", '-'), -- i=2177
      ("1001010001100111", '-'), -- i=2178
      ("1010010001100111", '-'), -- i=2179
      ("1011010001100111", '-'), -- i=2180
      ("0101010001100000", '1'), -- i=2181
      ("0100010001100000", '-'), -- i=2182
      ("0000010011101001", '-'), -- i=2183
      ("1000010001110000", '-'), -- i=2184
      ("1001010001110000", '-'), -- i=2185
      ("1010010001110000", '-'), -- i=2186
      ("1011010001110000", '-'), -- i=2187
      ("0101010001110000", '1'), -- i=2188
      ("0100010001110000", '-'), -- i=2189
      ("0000010011001010", '-'), -- i=2190
      ("1000010001110001", '-'), -- i=2191
      ("1001010001110001", '-'), -- i=2192
      ("1010010001110001", '-'), -- i=2193
      ("1011010001110001", '-'), -- i=2194
      ("0101010001110000", '1'), -- i=2195
      ("0100010001110000", '-'), -- i=2196
      ("0000010011100001", '-'), -- i=2197
      ("1000010001110010", '-'), -- i=2198
      ("1001010001110010", '-'), -- i=2199
      ("1010010001110010", '-'), -- i=2200
      ("1011010001110010", '-'), -- i=2201
      ("0101010001110000", '1'), -- i=2202
      ("0100010001110000", '-'), -- i=2203
      ("0000010001000001", '-'), -- i=2204
      ("1000010001110011", '-'), -- i=2205
      ("1001010001110011", '-'), -- i=2206
      ("1010010001110011", '-'), -- i=2207
      ("1011010001110011", '-'), -- i=2208
      ("0101010001110000", '1'), -- i=2209
      ("0100010001110000", '-'), -- i=2210
      ("0000010001101000", '-'), -- i=2211
      ("1000010001110100", '-'), -- i=2212
      ("1001010001110100", '-'), -- i=2213
      ("1010010001110100", '-'), -- i=2214
      ("1011010001110100", '-'), -- i=2215
      ("0101010001110000", '1'), -- i=2216
      ("0100010001110000", '-'), -- i=2217
      ("0000010011001110", '-'), -- i=2218
      ("1000010001110101", '-'), -- i=2219
      ("1001010001110101", '-'), -- i=2220
      ("1010010001110101", '-'), -- i=2221
      ("1011010001110101", '-'), -- i=2222
      ("0101010001110000", '1'), -- i=2223
      ("0100010001110000", '-'), -- i=2224
      ("0000010010001001", '-'), -- i=2225
      ("1000010001110110", '-'), -- i=2226
      ("1001010001110110", '-'), -- i=2227
      ("1010010001110110", '-'), -- i=2228
      ("1011010001110110", '-'), -- i=2229
      ("0101010001110000", '1'), -- i=2230
      ("0100010001110000", '-'), -- i=2231
      ("0000010010111001", '-'), -- i=2232
      ("1000010001110111", '-'), -- i=2233
      ("1001010001110111", '-'), -- i=2234
      ("1010010001110111", '-'), -- i=2235
      ("1011010001110111", '-'), -- i=2236
      ("0101010001110000", '1'), -- i=2237
      ("0100010001110000", '-'), -- i=2238
      ("0000010001111110", '-'), -- i=2239
      ("1000010100000000", '-'), -- i=2240
      ("1001010100000000", '-'), -- i=2241
      ("1010010100000000", '-'), -- i=2242
      ("1011010100000000", '-'), -- i=2243
      ("0101010100000000", '1'), -- i=2244
      ("0100010100000000", '-'), -- i=2245
      ("0000010111010000", '-'), -- i=2246
      ("1000010100000001", '-'), -- i=2247
      ("1001010100000001", '-'), -- i=2248
      ("1010010100000001", '-'), -- i=2249
      ("1011010100000001", '-'), -- i=2250
      ("0101010100000000", '1'), -- i=2251
      ("0100010100000000", '-'), -- i=2252
      ("0000010100110111", '-'), -- i=2253
      ("1000010100000010", '-'), -- i=2254
      ("1001010100000010", '-'), -- i=2255
      ("1010010100000010", '-'), -- i=2256
      ("1011010100000010", '-'), -- i=2257
      ("0101010100000000", '1'), -- i=2258
      ("0100010100000000", '-'), -- i=2259
      ("0000010101010100", '-'), -- i=2260
      ("1000010100000011", '-'), -- i=2261
      ("1001010100000011", '-'), -- i=2262
      ("1010010100000011", '-'), -- i=2263
      ("1011010100000011", '-'), -- i=2264
      ("0101010100000000", '1'), -- i=2265
      ("0100010100000000", '-'), -- i=2266
      ("0000010101110000", '-'), -- i=2267
      ("1000010100000100", '-'), -- i=2268
      ("1001010100000100", '-'), -- i=2269
      ("1010010100000100", '-'), -- i=2270
      ("1011010100000100", '-'), -- i=2271
      ("0101010100000000", '1'), -- i=2272
      ("0100010100000000", '-'), -- i=2273
      ("0000010111100000", '-'), -- i=2274
      ("1000010100000101", '-'), -- i=2275
      ("1001010100000101", '-'), -- i=2276
      ("1010010100000101", '-'), -- i=2277
      ("1011010100000101", '-'), -- i=2278
      ("0101010100000000", '1'), -- i=2279
      ("0100010100000000", '-'), -- i=2280
      ("0000010110100111", '-'), -- i=2281
      ("1000010100000110", '-'), -- i=2282
      ("1001010100000110", '-'), -- i=2283
      ("1010010100000110", '-'), -- i=2284
      ("1011010100000110", '-'), -- i=2285
      ("0101010100000000", '1'), -- i=2286
      ("0100010100000000", '-'), -- i=2287
      ("0000010111101111", '-'), -- i=2288
      ("1000010100000111", '-'), -- i=2289
      ("1001010100000111", '-'), -- i=2290
      ("1010010100000111", '-'), -- i=2291
      ("1011010100000111", '-'), -- i=2292
      ("0101010100000000", '1'), -- i=2293
      ("0100010100000000", '-'), -- i=2294
      ("0000010101110000", '-'), -- i=2295
      ("1000010100010000", '-'), -- i=2296
      ("1001010100010000", '-'), -- i=2297
      ("1010010100010000", '-'), -- i=2298
      ("1011010100010000", '-'), -- i=2299
      ("0101010100010000", '1'), -- i=2300
      ("0100010100010000", '-'), -- i=2301
      ("0000010111111011", '-'), -- i=2302
      ("1000010100010001", '-'), -- i=2303
      ("1001010100010001", '-'), -- i=2304
      ("1010010100010001", '-'), -- i=2305
      ("1011010100010001", '-'), -- i=2306
      ("0101010100010000", '1'), -- i=2307
      ("0100010100010000", '-'), -- i=2308
      ("0000010111101100", '-'), -- i=2309
      ("1000010100010010", '-'), -- i=2310
      ("1001010100010010", '-'), -- i=2311
      ("1010010100010010", '-'), -- i=2312
      ("1011010100010010", '-'), -- i=2313
      ("0101010100010000", '1'), -- i=2314
      ("0100010100010000", '-'), -- i=2315
      ("0000010111100011", '-'), -- i=2316
      ("1000010100010011", '-'), -- i=2317
      ("1001010100010011", '-'), -- i=2318
      ("1010010100010011", '-'), -- i=2319
      ("1011010100010011", '-'), -- i=2320
      ("0101010100010000", '1'), -- i=2321
      ("0100010100010000", '-'), -- i=2322
      ("0000010110001101", '-'), -- i=2323
      ("1000010100010100", '-'), -- i=2324
      ("1001010100010100", '-'), -- i=2325
      ("1010010100010100", '-'), -- i=2326
      ("1011010100010100", '-'), -- i=2327
      ("0101010100010000", '1'), -- i=2328
      ("0100010100010000", '-'), -- i=2329
      ("0000010111010111", '-'), -- i=2330
      ("1000010100010101", '-'), -- i=2331
      ("1001010100010101", '-'), -- i=2332
      ("1010010100010101", '-'), -- i=2333
      ("1011010100010101", '-'), -- i=2334
      ("0101010100010000", '1'), -- i=2335
      ("0100010100010000", '-'), -- i=2336
      ("0000010100101010", '-'), -- i=2337
      ("1000010100010110", '-'), -- i=2338
      ("1001010100010110", '-'), -- i=2339
      ("1010010100010110", '-'), -- i=2340
      ("1011010100010110", '-'), -- i=2341
      ("0101010100010000", '1'), -- i=2342
      ("0100010100010000", '-'), -- i=2343
      ("0000010110011110", '-'), -- i=2344
      ("1000010100010111", '-'), -- i=2345
      ("1001010100010111", '-'), -- i=2346
      ("1010010100010111", '-'), -- i=2347
      ("1011010100010111", '-'), -- i=2348
      ("0101010100010000", '1'), -- i=2349
      ("0100010100010000", '-'), -- i=2350
      ("0000010100011100", '-'), -- i=2351
      ("1000010100100000", '-'), -- i=2352
      ("1001010100100000", '-'), -- i=2353
      ("1010010100100000", '-'), -- i=2354
      ("1011010100100000", '-'), -- i=2355
      ("0101010100100000", '1'), -- i=2356
      ("0100010100100000", '-'), -- i=2357
      ("0000010110110101", '-'), -- i=2358
      ("1000010100100001", '-'), -- i=2359
      ("1001010100100001", '-'), -- i=2360
      ("1010010100100001", '-'), -- i=2361
      ("1011010100100001", '-'), -- i=2362
      ("0101010100100000", '1'), -- i=2363
      ("0100010100100000", '-'), -- i=2364
      ("0000010100100111", '-'), -- i=2365
      ("1000010100100010", '-'), -- i=2366
      ("1001010100100010", '-'), -- i=2367
      ("1010010100100010", '-'), -- i=2368
      ("1011010100100010", '-'), -- i=2369
      ("0101010100100000", '1'), -- i=2370
      ("0100010100100000", '-'), -- i=2371
      ("0000010101111010", '-'), -- i=2372
      ("1000010100100011", '-'), -- i=2373
      ("1001010100100011", '-'), -- i=2374
      ("1010010100100011", '-'), -- i=2375
      ("1011010100100011", '-'), -- i=2376
      ("0101010100100000", '1'), -- i=2377
      ("0100010100100000", '-'), -- i=2378
      ("0000010110000111", '-'), -- i=2379
      ("1000010100100100", '-'), -- i=2380
      ("1001010100100100", '-'), -- i=2381
      ("1010010100100100", '-'), -- i=2382
      ("1011010100100100", '-'), -- i=2383
      ("0101010100100000", '1'), -- i=2384
      ("0100010100100000", '-'), -- i=2385
      ("0000010101011101", '-'), -- i=2386
      ("1000010100100101", '-'), -- i=2387
      ("1001010100100101", '-'), -- i=2388
      ("1010010100100101", '-'), -- i=2389
      ("1011010100100101", '-'), -- i=2390
      ("0101010100100000", '1'), -- i=2391
      ("0100010100100000", '-'), -- i=2392
      ("0000010100011011", '-'), -- i=2393
      ("1000010100100110", '-'), -- i=2394
      ("1001010100100110", '-'), -- i=2395
      ("1010010100100110", '-'), -- i=2396
      ("1011010100100110", '-'), -- i=2397
      ("0101010100100000", '1'), -- i=2398
      ("0100010100100000", '-'), -- i=2399
      ("0000010101011010", '-'), -- i=2400
      ("1000010100100111", '-'), -- i=2401
      ("1001010100100111", '-'), -- i=2402
      ("1010010100100111", '-'), -- i=2403
      ("1011010100100111", '-'), -- i=2404
      ("0101010100100000", '1'), -- i=2405
      ("0100010100100000", '-'), -- i=2406
      ("0000010111000111", '-'), -- i=2407
      ("1000010100110000", '-'), -- i=2408
      ("1001010100110000", '-'), -- i=2409
      ("1010010100110000", '-'), -- i=2410
      ("1011010100110000", '-'), -- i=2411
      ("0101010100110000", '1'), -- i=2412
      ("0100010100110000", '-'), -- i=2413
      ("0000010111000101", '-'), -- i=2414
      ("1000010100110001", '-'), -- i=2415
      ("1001010100110001", '-'), -- i=2416
      ("1010010100110001", '-'), -- i=2417
      ("1011010100110001", '-'), -- i=2418
      ("0101010100110000", '1'), -- i=2419
      ("0100010100110000", '-'), -- i=2420
      ("0000010100110100", '-'), -- i=2421
      ("1000010100110010", '-'), -- i=2422
      ("1001010100110010", '-'), -- i=2423
      ("1010010100110010", '-'), -- i=2424
      ("1011010100110010", '-'), -- i=2425
      ("0101010100110000", '1'), -- i=2426
      ("0100010100110000", '-'), -- i=2427
      ("0000010100100110", '-'), -- i=2428
      ("1000010100110011", '-'), -- i=2429
      ("1001010100110011", '-'), -- i=2430
      ("1010010100110011", '-'), -- i=2431
      ("1011010100110011", '-'), -- i=2432
      ("0101010100110000", '1'), -- i=2433
      ("0100010100110000", '-'), -- i=2434
      ("0000010101011111", '-'), -- i=2435
      ("1000010100110100", '-'), -- i=2436
      ("1001010100110100", '-'), -- i=2437
      ("1010010100110100", '-'), -- i=2438
      ("1011010100110100", '-'), -- i=2439
      ("0101010100110000", '1'), -- i=2440
      ("0100010100110000", '-'), -- i=2441
      ("0000010110101111", '-'), -- i=2442
      ("1000010100110101", '-'), -- i=2443
      ("1001010100110101", '-'), -- i=2444
      ("1010010100110101", '-'), -- i=2445
      ("1011010100110101", '-'), -- i=2446
      ("0101010100110000", '1'), -- i=2447
      ("0100010100110000", '-'), -- i=2448
      ("0000010110110000", '-'), -- i=2449
      ("1000010100110110", '-'), -- i=2450
      ("1001010100110110", '-'), -- i=2451
      ("1010010100110110", '-'), -- i=2452
      ("1011010100110110", '-'), -- i=2453
      ("0101010100110000", '1'), -- i=2454
      ("0100010100110000", '-'), -- i=2455
      ("0000010110100000", '-'), -- i=2456
      ("1000010100110111", '-'), -- i=2457
      ("1001010100110111", '-'), -- i=2458
      ("1010010100110111", '-'), -- i=2459
      ("1011010100110111", '-'), -- i=2460
      ("0101010100110000", '1'), -- i=2461
      ("0100010100110000", '-'), -- i=2462
      ("0000010110111001", '-'), -- i=2463
      ("1000010101000000", '-'), -- i=2464
      ("1001010101000000", '-'), -- i=2465
      ("1010010101000000", '-'), -- i=2466
      ("1011010101000000", '-'), -- i=2467
      ("0101010101000000", '1'), -- i=2468
      ("0100010101000000", '-'), -- i=2469
      ("0000010100011100", '-'), -- i=2470
      ("1000010101000001", '-'), -- i=2471
      ("1001010101000001", '-'), -- i=2472
      ("1010010101000001", '-'), -- i=2473
      ("1011010101000001", '-'), -- i=2474
      ("0101010101000000", '1'), -- i=2475
      ("0100010101000000", '-'), -- i=2476
      ("0000010100100000", '-'), -- i=2477
      ("1000010101000010", '-'), -- i=2478
      ("1001010101000010", '-'), -- i=2479
      ("1010010101000010", '-'), -- i=2480
      ("1011010101000010", '-'), -- i=2481
      ("0101010101000000", '1'), -- i=2482
      ("0100010101000000", '-'), -- i=2483
      ("0000010111000001", '-'), -- i=2484
      ("1000010101000011", '-'), -- i=2485
      ("1001010101000011", '-'), -- i=2486
      ("1010010101000011", '-'), -- i=2487
      ("1011010101000011", '-'), -- i=2488
      ("0101010101000000", '1'), -- i=2489
      ("0100010101000000", '-'), -- i=2490
      ("0000010111011110", '-'), -- i=2491
      ("1000010101000100", '-'), -- i=2492
      ("1001010101000100", '-'), -- i=2493
      ("1010010101000100", '-'), -- i=2494
      ("1011010101000100", '-'), -- i=2495
      ("0101010101000000", '1'), -- i=2496
      ("0100010101000000", '-'), -- i=2497
      ("0000010100100111", '-'), -- i=2498
      ("1000010101000101", '-'), -- i=2499
      ("1001010101000101", '-'), -- i=2500
      ("1010010101000101", '-'), -- i=2501
      ("1011010101000101", '-'), -- i=2502
      ("0101010101000000", '1'), -- i=2503
      ("0100010101000000", '-'), -- i=2504
      ("0000010101011111", '-'), -- i=2505
      ("1000010101000110", '-'), -- i=2506
      ("1001010101000110", '-'), -- i=2507
      ("1010010101000110", '-'), -- i=2508
      ("1011010101000110", '-'), -- i=2509
      ("0101010101000000", '1'), -- i=2510
      ("0100010101000000", '-'), -- i=2511
      ("0000010100110111", '-'), -- i=2512
      ("1000010101000111", '-'), -- i=2513
      ("1001010101000111", '-'), -- i=2514
      ("1010010101000111", '-'), -- i=2515
      ("1011010101000111", '-'), -- i=2516
      ("0101010101000000", '1'), -- i=2517
      ("0100010101000000", '-'), -- i=2518
      ("0000010100011011", '-'), -- i=2519
      ("1000010101010000", '-'), -- i=2520
      ("1001010101010000", '-'), -- i=2521
      ("1010010101010000", '-'), -- i=2522
      ("1011010101010000", '-'), -- i=2523
      ("0101010101010000", '1'), -- i=2524
      ("0100010101010000", '-'), -- i=2525
      ("0000010101111101", '-'), -- i=2526
      ("1000010101010001", '-'), -- i=2527
      ("1001010101010001", '-'), -- i=2528
      ("1010010101010001", '-'), -- i=2529
      ("1011010101010001", '-'), -- i=2530
      ("0101010101010000", '1'), -- i=2531
      ("0100010101010000", '-'), -- i=2532
      ("0000010100000111", '-'), -- i=2533
      ("1000010101010010", '-'), -- i=2534
      ("1001010101010010", '-'), -- i=2535
      ("1010010101010010", '-'), -- i=2536
      ("1011010101010010", '-'), -- i=2537
      ("0101010101010000", '1'), -- i=2538
      ("0100010101010000", '-'), -- i=2539
      ("0000010101000100", '-'), -- i=2540
      ("1000010101010011", '-'), -- i=2541
      ("1001010101010011", '-'), -- i=2542
      ("1010010101010011", '-'), -- i=2543
      ("1011010101010011", '-'), -- i=2544
      ("0101010101010000", '1'), -- i=2545
      ("0100010101010000", '-'), -- i=2546
      ("0000010110111111", '-'), -- i=2547
      ("1000010101010100", '-'), -- i=2548
      ("1001010101010100", '-'), -- i=2549
      ("1010010101010100", '-'), -- i=2550
      ("1011010101010100", '-'), -- i=2551
      ("0101010101010000", '1'), -- i=2552
      ("0100010101010000", '-'), -- i=2553
      ("0000010110010011", '-'), -- i=2554
      ("1000010101010101", '-'), -- i=2555
      ("1001010101010101", '-'), -- i=2556
      ("1010010101010101", '-'), -- i=2557
      ("1011010101010101", '-'), -- i=2558
      ("0101010101010000", '1'), -- i=2559
      ("0100010101010000", '-'), -- i=2560
      ("0000010110111001", '-'), -- i=2561
      ("1000010101010110", '-'), -- i=2562
      ("1001010101010110", '-'), -- i=2563
      ("1010010101010110", '-'), -- i=2564
      ("1011010101010110", '-'), -- i=2565
      ("0101010101010000", '1'), -- i=2566
      ("0100010101010000", '-'), -- i=2567
      ("0000010111111110", '-'), -- i=2568
      ("1000010101010111", '-'), -- i=2569
      ("1001010101010111", '-'), -- i=2570
      ("1010010101010111", '-'), -- i=2571
      ("1011010101010111", '-'), -- i=2572
      ("0101010101010000", '1'), -- i=2573
      ("0100010101010000", '-'), -- i=2574
      ("0000010101011111", '-'), -- i=2575
      ("1000010101100000", '-'), -- i=2576
      ("1001010101100000", '-'), -- i=2577
      ("1010010101100000", '-'), -- i=2578
      ("1011010101100000", '-'), -- i=2579
      ("0101010101100000", '1'), -- i=2580
      ("0100010101100000", '-'), -- i=2581
      ("0000010101001011", '-'), -- i=2582
      ("1000010101100001", '-'), -- i=2583
      ("1001010101100001", '-'), -- i=2584
      ("1010010101100001", '-'), -- i=2585
      ("1011010101100001", '-'), -- i=2586
      ("0101010101100000", '1'), -- i=2587
      ("0100010101100000", '-'), -- i=2588
      ("0000010101010010", '-'), -- i=2589
      ("1000010101100010", '-'), -- i=2590
      ("1001010101100010", '-'), -- i=2591
      ("1010010101100010", '-'), -- i=2592
      ("1011010101100010", '-'), -- i=2593
      ("0101010101100000", '1'), -- i=2594
      ("0100010101100000", '-'), -- i=2595
      ("0000010101100010", '-'), -- i=2596
      ("1000010101100011", '-'), -- i=2597
      ("1001010101100011", '-'), -- i=2598
      ("1010010101100011", '-'), -- i=2599
      ("1011010101100011", '-'), -- i=2600
      ("0101010101100000", '1'), -- i=2601
      ("0100010101100000", '-'), -- i=2602
      ("0000010100111000", '-'), -- i=2603
      ("1000010101100100", '-'), -- i=2604
      ("1001010101100100", '-'), -- i=2605
      ("1010010101100100", '-'), -- i=2606
      ("1011010101100100", '-'), -- i=2607
      ("0101010101100000", '1'), -- i=2608
      ("0100010101100000", '-'), -- i=2609
      ("0000010110101110", '-'), -- i=2610
      ("1000010101100101", '-'), -- i=2611
      ("1001010101100101", '-'), -- i=2612
      ("1010010101100101", '-'), -- i=2613
      ("1011010101100101", '-'), -- i=2614
      ("0101010101100000", '1'), -- i=2615
      ("0100010101100000", '-'), -- i=2616
      ("0000010101100011", '-'), -- i=2617
      ("1000010101100110", '-'), -- i=2618
      ("1001010101100110", '-'), -- i=2619
      ("1010010101100110", '-'), -- i=2620
      ("1011010101100110", '-'), -- i=2621
      ("0101010101100000", '1'), -- i=2622
      ("0100010101100000", '-'), -- i=2623
      ("0000010110010011", '-'), -- i=2624
      ("1000010101100111", '-'), -- i=2625
      ("1001010101100111", '-'), -- i=2626
      ("1010010101100111", '-'), -- i=2627
      ("1011010101100111", '-'), -- i=2628
      ("0101010101100000", '1'), -- i=2629
      ("0100010101100000", '-'), -- i=2630
      ("0000010111110101", '-'), -- i=2631
      ("1000010101110000", '-'), -- i=2632
      ("1001010101110000", '-'), -- i=2633
      ("1010010101110000", '-'), -- i=2634
      ("1011010101110000", '-'), -- i=2635
      ("0101010101110000", '1'), -- i=2636
      ("0100010101110000", '-'), -- i=2637
      ("0000010100100011", '-'), -- i=2638
      ("1000010101110001", '-'), -- i=2639
      ("1001010101110001", '-'), -- i=2640
      ("1010010101110001", '-'), -- i=2641
      ("1011010101110001", '-'), -- i=2642
      ("0101010101110000", '1'), -- i=2643
      ("0100010101110000", '-'), -- i=2644
      ("0000010101010111", '-'), -- i=2645
      ("1000010101110010", '-'), -- i=2646
      ("1001010101110010", '-'), -- i=2647
      ("1010010101110010", '-'), -- i=2648
      ("1011010101110010", '-'), -- i=2649
      ("0101010101110000", '1'), -- i=2650
      ("0100010101110000", '-'), -- i=2651
      ("0000010100110011", '-'), -- i=2652
      ("1000010101110011", '-'), -- i=2653
      ("1001010101110011", '-'), -- i=2654
      ("1010010101110011", '-'), -- i=2655
      ("1011010101110011", '-'), -- i=2656
      ("0101010101110000", '1'), -- i=2657
      ("0100010101110000", '-'), -- i=2658
      ("0000010111111011", '-'), -- i=2659
      ("1000010101110100", '-'), -- i=2660
      ("1001010101110100", '-'), -- i=2661
      ("1010010101110100", '-'), -- i=2662
      ("1011010101110100", '-'), -- i=2663
      ("0101010101110000", '1'), -- i=2664
      ("0100010101110000", '-'), -- i=2665
      ("0000010101111100", '-'), -- i=2666
      ("1000010101110101", '-'), -- i=2667
      ("1001010101110101", '-'), -- i=2668
      ("1010010101110101", '-'), -- i=2669
      ("1011010101110101", '-'), -- i=2670
      ("0101010101110000", '1'), -- i=2671
      ("0100010101110000", '-'), -- i=2672
      ("0000010111001101", '-'), -- i=2673
      ("1000010101110110", '-'), -- i=2674
      ("1001010101110110", '-'), -- i=2675
      ("1010010101110110", '-'), -- i=2676
      ("1011010101110110", '-'), -- i=2677
      ("0101010101110000", '1'), -- i=2678
      ("0100010101110000", '-'), -- i=2679
      ("0000010110100101", '-'), -- i=2680
      ("1000010101110111", '-'), -- i=2681
      ("1001010101110111", '-'), -- i=2682
      ("1010010101110111", '-'), -- i=2683
      ("1011010101110111", '-'), -- i=2684
      ("0101010101110000", '1'), -- i=2685
      ("0100010101110000", '-'), -- i=2686
      ("0000010110011010", '-'), -- i=2687
      ("1000011000000000", '-'), -- i=2688
      ("1001011000000000", '-'), -- i=2689
      ("1010011000000000", '-'), -- i=2690
      ("1011011000000000", '-'), -- i=2691
      ("0101011000000000", '1'), -- i=2692
      ("0100011000000000", '-'), -- i=2693
      ("0000011011111000", '-'), -- i=2694
      ("1000011000000001", '-'), -- i=2695
      ("1001011000000001", '-'), -- i=2696
      ("1010011000000001", '-'), -- i=2697
      ("1011011000000001", '-'), -- i=2698
      ("0101011000000000", '1'), -- i=2699
      ("0100011000000000", '-'), -- i=2700
      ("0000011000010101", '-'), -- i=2701
      ("1000011000000010", '-'), -- i=2702
      ("1001011000000010", '-'), -- i=2703
      ("1010011000000010", '-'), -- i=2704
      ("1011011000000010", '-'), -- i=2705
      ("0101011000000000", '1'), -- i=2706
      ("0100011000000000", '-'), -- i=2707
      ("0000011010101111", '-'), -- i=2708
      ("1000011000000011", '-'), -- i=2709
      ("1001011000000011", '-'), -- i=2710
      ("1010011000000011", '-'), -- i=2711
      ("1011011000000011", '-'), -- i=2712
      ("0101011000000000", '1'), -- i=2713
      ("0100011000000000", '-'), -- i=2714
      ("0000011011011110", '-'), -- i=2715
      ("1000011000000100", '-'), -- i=2716
      ("1001011000000100", '-'), -- i=2717
      ("1010011000000100", '-'), -- i=2718
      ("1011011000000100", '-'), -- i=2719
      ("0101011000000000", '1'), -- i=2720
      ("0100011000000000", '-'), -- i=2721
      ("0000011001110110", '-'), -- i=2722
      ("1000011000000101", '-'), -- i=2723
      ("1001011000000101", '-'), -- i=2724
      ("1010011000000101", '-'), -- i=2725
      ("1011011000000101", '-'), -- i=2726
      ("0101011000000000", '1'), -- i=2727
      ("0100011000000000", '-'), -- i=2728
      ("0000011001110111", '-'), -- i=2729
      ("1000011000000110", '-'), -- i=2730
      ("1001011000000110", '-'), -- i=2731
      ("1010011000000110", '-'), -- i=2732
      ("1011011000000110", '-'), -- i=2733
      ("0101011000000000", '1'), -- i=2734
      ("0100011000000000", '-'), -- i=2735
      ("0000011011101100", '-'), -- i=2736
      ("1000011000000111", '-'), -- i=2737
      ("1001011000000111", '-'), -- i=2738
      ("1010011000000111", '-'), -- i=2739
      ("1011011000000111", '-'), -- i=2740
      ("0101011000000000", '1'), -- i=2741
      ("0100011000000000", '-'), -- i=2742
      ("0000011010001110", '-'), -- i=2743
      ("1000011000010000", '-'), -- i=2744
      ("1001011000010000", '-'), -- i=2745
      ("1010011000010000", '-'), -- i=2746
      ("1011011000010000", '-'), -- i=2747
      ("0101011000010000", '1'), -- i=2748
      ("0100011000010000", '-'), -- i=2749
      ("0000011011010111", '-'), -- i=2750
      ("1000011000010001", '-'), -- i=2751
      ("1001011000010001", '-'), -- i=2752
      ("1010011000010001", '-'), -- i=2753
      ("1011011000010001", '-'), -- i=2754
      ("0101011000010000", '1'), -- i=2755
      ("0100011000010000", '-'), -- i=2756
      ("0000011000001010", '-'), -- i=2757
      ("1000011000010010", '-'), -- i=2758
      ("1001011000010010", '-'), -- i=2759
      ("1010011000010010", '-'), -- i=2760
      ("1011011000010010", '-'), -- i=2761
      ("0101011000010000", '1'), -- i=2762
      ("0100011000010000", '-'), -- i=2763
      ("0000011000101110", '-'), -- i=2764
      ("1000011000010011", '-'), -- i=2765
      ("1001011000010011", '-'), -- i=2766
      ("1010011000010011", '-'), -- i=2767
      ("1011011000010011", '-'), -- i=2768
      ("0101011000010000", '1'), -- i=2769
      ("0100011000010000", '-'), -- i=2770
      ("0000011011010010", '-'), -- i=2771
      ("1000011000010100", '-'), -- i=2772
      ("1001011000010100", '-'), -- i=2773
      ("1010011000010100", '-'), -- i=2774
      ("1011011000010100", '-'), -- i=2775
      ("0101011000010000", '1'), -- i=2776
      ("0100011000010000", '-'), -- i=2777
      ("0000011010111001", '-'), -- i=2778
      ("1000011000010101", '-'), -- i=2779
      ("1001011000010101", '-'), -- i=2780
      ("1010011000010101", '-'), -- i=2781
      ("1011011000010101", '-'), -- i=2782
      ("0101011000010000", '1'), -- i=2783
      ("0100011000010000", '-'), -- i=2784
      ("0000011011100011", '-'), -- i=2785
      ("1000011000010110", '-'), -- i=2786
      ("1001011000010110", '-'), -- i=2787
      ("1010011000010110", '-'), -- i=2788
      ("1011011000010110", '-'), -- i=2789
      ("0101011000010000", '1'), -- i=2790
      ("0100011000010000", '-'), -- i=2791
      ("0000011000000011", '-'), -- i=2792
      ("1000011000010111", '-'), -- i=2793
      ("1001011000010111", '-'), -- i=2794
      ("1010011000010111", '-'), -- i=2795
      ("1011011000010111", '-'), -- i=2796
      ("0101011000010000", '1'), -- i=2797
      ("0100011000010000", '-'), -- i=2798
      ("0000011001101100", '-'), -- i=2799
      ("1000011000100000", '-'), -- i=2800
      ("1001011000100000", '-'), -- i=2801
      ("1010011000100000", '-'), -- i=2802
      ("1011011000100000", '-'), -- i=2803
      ("0101011000100000", '1'), -- i=2804
      ("0100011000100000", '-'), -- i=2805
      ("0000011010011010", '-'), -- i=2806
      ("1000011000100001", '-'), -- i=2807
      ("1001011000100001", '-'), -- i=2808
      ("1010011000100001", '-'), -- i=2809
      ("1011011000100001", '-'), -- i=2810
      ("0101011000100000", '1'), -- i=2811
      ("0100011000100000", '-'), -- i=2812
      ("0000011001011010", '-'), -- i=2813
      ("1000011000100010", '-'), -- i=2814
      ("1001011000100010", '-'), -- i=2815
      ("1010011000100010", '-'), -- i=2816
      ("1011011000100010", '-'), -- i=2817
      ("0101011000100000", '1'), -- i=2818
      ("0100011000100000", '-'), -- i=2819
      ("0000011001000011", '-'), -- i=2820
      ("1000011000100011", '-'), -- i=2821
      ("1001011000100011", '-'), -- i=2822
      ("1010011000100011", '-'), -- i=2823
      ("1011011000100011", '-'), -- i=2824
      ("0101011000100000", '1'), -- i=2825
      ("0100011000100000", '-'), -- i=2826
      ("0000011011010011", '-'), -- i=2827
      ("1000011000100100", '-'), -- i=2828
      ("1001011000100100", '-'), -- i=2829
      ("1010011000100100", '-'), -- i=2830
      ("1011011000100100", '-'), -- i=2831
      ("0101011000100000", '1'), -- i=2832
      ("0100011000100000", '-'), -- i=2833
      ("0000011010011110", '-'), -- i=2834
      ("1000011000100101", '-'), -- i=2835
      ("1001011000100101", '-'), -- i=2836
      ("1010011000100101", '-'), -- i=2837
      ("1011011000100101", '-'), -- i=2838
      ("0101011000100000", '1'), -- i=2839
      ("0100011000100000", '-'), -- i=2840
      ("0000011010001010", '-'), -- i=2841
      ("1000011000100110", '-'), -- i=2842
      ("1001011000100110", '-'), -- i=2843
      ("1010011000100110", '-'), -- i=2844
      ("1011011000100110", '-'), -- i=2845
      ("0101011000100000", '1'), -- i=2846
      ("0100011000100000", '-'), -- i=2847
      ("0000011010110010", '-'), -- i=2848
      ("1000011000100111", '-'), -- i=2849
      ("1001011000100111", '-'), -- i=2850
      ("1010011000100111", '-'), -- i=2851
      ("1011011000100111", '-'), -- i=2852
      ("0101011000100000", '1'), -- i=2853
      ("0100011000100000", '-'), -- i=2854
      ("0000011010000100", '-'), -- i=2855
      ("1000011000110000", '-'), -- i=2856
      ("1001011000110000", '-'), -- i=2857
      ("1010011000110000", '-'), -- i=2858
      ("1011011000110000", '-'), -- i=2859
      ("0101011000110000", '1'), -- i=2860
      ("0100011000110000", '-'), -- i=2861
      ("0000011000011101", '-'), -- i=2862
      ("1000011000110001", '-'), -- i=2863
      ("1001011000110001", '-'), -- i=2864
      ("1010011000110001", '-'), -- i=2865
      ("1011011000110001", '-'), -- i=2866
      ("0101011000110000", '1'), -- i=2867
      ("0100011000110000", '-'), -- i=2868
      ("0000011010111001", '-'), -- i=2869
      ("1000011000110010", '-'), -- i=2870
      ("1001011000110010", '-'), -- i=2871
      ("1010011000110010", '-'), -- i=2872
      ("1011011000110010", '-'), -- i=2873
      ("0101011000110000", '1'), -- i=2874
      ("0100011000110000", '-'), -- i=2875
      ("0000011010011010", '-'), -- i=2876
      ("1000011000110011", '-'), -- i=2877
      ("1001011000110011", '-'), -- i=2878
      ("1010011000110011", '-'), -- i=2879
      ("1011011000110011", '-'), -- i=2880
      ("0101011000110000", '1'), -- i=2881
      ("0100011000110000", '-'), -- i=2882
      ("0000011011110100", '-'), -- i=2883
      ("1000011000110100", '-'), -- i=2884
      ("1001011000110100", '-'), -- i=2885
      ("1010011000110100", '-'), -- i=2886
      ("1011011000110100", '-'), -- i=2887
      ("0101011000110000", '1'), -- i=2888
      ("0100011000110000", '-'), -- i=2889
      ("0000011001111111", '-'), -- i=2890
      ("1000011000110101", '-'), -- i=2891
      ("1001011000110101", '-'), -- i=2892
      ("1010011000110101", '-'), -- i=2893
      ("1011011000110101", '-'), -- i=2894
      ("0101011000110000", '1'), -- i=2895
      ("0100011000110000", '-'), -- i=2896
      ("0000011001101111", '-'), -- i=2897
      ("1000011000110110", '-'), -- i=2898
      ("1001011000110110", '-'), -- i=2899
      ("1010011000110110", '-'), -- i=2900
      ("1011011000110110", '-'), -- i=2901
      ("0101011000110000", '1'), -- i=2902
      ("0100011000110000", '-'), -- i=2903
      ("0000011001010110", '-'), -- i=2904
      ("1000011000110111", '-'), -- i=2905
      ("1001011000110111", '-'), -- i=2906
      ("1010011000110111", '-'), -- i=2907
      ("1011011000110111", '-'), -- i=2908
      ("0101011000110000", '1'), -- i=2909
      ("0100011000110000", '-'), -- i=2910
      ("0000011011100011", '-'), -- i=2911
      ("1000011001000000", '-'), -- i=2912
      ("1001011001000000", '-'), -- i=2913
      ("1010011001000000", '-'), -- i=2914
      ("1011011001000000", '-'), -- i=2915
      ("0101011001000000", '1'), -- i=2916
      ("0100011001000000", '-'), -- i=2917
      ("0000011011000011", '-'), -- i=2918
      ("1000011001000001", '-'), -- i=2919
      ("1001011001000001", '-'), -- i=2920
      ("1010011001000001", '-'), -- i=2921
      ("1011011001000001", '-'), -- i=2922
      ("0101011001000000", '1'), -- i=2923
      ("0100011001000000", '-'), -- i=2924
      ("0000011011011110", '-'), -- i=2925
      ("1000011001000010", '-'), -- i=2926
      ("1001011001000010", '-'), -- i=2927
      ("1010011001000010", '-'), -- i=2928
      ("1011011001000010", '-'), -- i=2929
      ("0101011001000000", '1'), -- i=2930
      ("0100011001000000", '-'), -- i=2931
      ("0000011010111011", '-'), -- i=2932
      ("1000011001000011", '-'), -- i=2933
      ("1001011001000011", '-'), -- i=2934
      ("1010011001000011", '-'), -- i=2935
      ("1011011001000011", '-'), -- i=2936
      ("0101011001000000", '1'), -- i=2937
      ("0100011001000000", '-'), -- i=2938
      ("0000011010111111", '-'), -- i=2939
      ("1000011001000100", '-'), -- i=2940
      ("1001011001000100", '-'), -- i=2941
      ("1010011001000100", '-'), -- i=2942
      ("1011011001000100", '-'), -- i=2943
      ("0101011001000000", '1'), -- i=2944
      ("0100011001000000", '-'), -- i=2945
      ("0000011010001001", '-'), -- i=2946
      ("1000011001000101", '-'), -- i=2947
      ("1001011001000101", '-'), -- i=2948
      ("1010011001000101", '-'), -- i=2949
      ("1011011001000101", '-'), -- i=2950
      ("0101011001000000", '1'), -- i=2951
      ("0100011001000000", '-'), -- i=2952
      ("0000011000101010", '-'), -- i=2953
      ("1000011001000110", '-'), -- i=2954
      ("1001011001000110", '-'), -- i=2955
      ("1010011001000110", '-'), -- i=2956
      ("1011011001000110", '-'), -- i=2957
      ("0101011001000000", '1'), -- i=2958
      ("0100011001000000", '-'), -- i=2959
      ("0000011010000000", '-'), -- i=2960
      ("1000011001000111", '-'), -- i=2961
      ("1001011001000111", '-'), -- i=2962
      ("1010011001000111", '-'), -- i=2963
      ("1011011001000111", '-'), -- i=2964
      ("0101011001000000", '1'), -- i=2965
      ("0100011001000000", '-'), -- i=2966
      ("0000011001110001", '-'), -- i=2967
      ("1000011001010000", '-'), -- i=2968
      ("1001011001010000", '-'), -- i=2969
      ("1010011001010000", '-'), -- i=2970
      ("1011011001010000", '-'), -- i=2971
      ("0101011001010000", '1'), -- i=2972
      ("0100011001010000", '-'), -- i=2973
      ("0000011001101000", '-'), -- i=2974
      ("1000011001010001", '-'), -- i=2975
      ("1001011001010001", '-'), -- i=2976
      ("1010011001010001", '-'), -- i=2977
      ("1011011001010001", '-'), -- i=2978
      ("0101011001010000", '1'), -- i=2979
      ("0100011001010000", '-'), -- i=2980
      ("0000011001100110", '-'), -- i=2981
      ("1000011001010010", '-'), -- i=2982
      ("1001011001010010", '-'), -- i=2983
      ("1010011001010010", '-'), -- i=2984
      ("1011011001010010", '-'), -- i=2985
      ("0101011001010000", '1'), -- i=2986
      ("0100011001010000", '-'), -- i=2987
      ("0000011011000100", '-'), -- i=2988
      ("1000011001010011", '-'), -- i=2989
      ("1001011001010011", '-'), -- i=2990
      ("1010011001010011", '-'), -- i=2991
      ("1011011001010011", '-'), -- i=2992
      ("0101011001010000", '1'), -- i=2993
      ("0100011001010000", '-'), -- i=2994
      ("0000011001111110", '-'), -- i=2995
      ("1000011001010100", '-'), -- i=2996
      ("1001011001010100", '-'), -- i=2997
      ("1010011001010100", '-'), -- i=2998
      ("1011011001010100", '-'), -- i=2999
      ("0101011001010000", '1'), -- i=3000
      ("0100011001010000", '-'), -- i=3001
      ("0000011011010111", '-'), -- i=3002
      ("1000011001010101", '-'), -- i=3003
      ("1001011001010101", '-'), -- i=3004
      ("1010011001010101", '-'), -- i=3005
      ("1011011001010101", '-'), -- i=3006
      ("0101011001010000", '1'), -- i=3007
      ("0100011001010000", '-'), -- i=3008
      ("0000011010000010", '-'), -- i=3009
      ("1000011001010110", '-'), -- i=3010
      ("1001011001010110", '-'), -- i=3011
      ("1010011001010110", '-'), -- i=3012
      ("1011011001010110", '-'), -- i=3013
      ("0101011001010000", '1'), -- i=3014
      ("0100011001010000", '-'), -- i=3015
      ("0000011011110011", '-'), -- i=3016
      ("1000011001010111", '-'), -- i=3017
      ("1001011001010111", '-'), -- i=3018
      ("1010011001010111", '-'), -- i=3019
      ("1011011001010111", '-'), -- i=3020
      ("0101011001010000", '1'), -- i=3021
      ("0100011001010000", '-'), -- i=3022
      ("0000011011001101", '-'), -- i=3023
      ("1000011001100000", '-'), -- i=3024
      ("1001011001100000", '-'), -- i=3025
      ("1010011001100000", '-'), -- i=3026
      ("1011011001100000", '-'), -- i=3027
      ("0101011001100000", '1'), -- i=3028
      ("0100011001100000", '-'), -- i=3029
      ("0000011011111100", '-'), -- i=3030
      ("1000011001100001", '-'), -- i=3031
      ("1001011001100001", '-'), -- i=3032
      ("1010011001100001", '-'), -- i=3033
      ("1011011001100001", '-'), -- i=3034
      ("0101011001100000", '1'), -- i=3035
      ("0100011001100000", '-'), -- i=3036
      ("0000011001111100", '-'), -- i=3037
      ("1000011001100010", '-'), -- i=3038
      ("1001011001100010", '-'), -- i=3039
      ("1010011001100010", '-'), -- i=3040
      ("1011011001100010", '-'), -- i=3041
      ("0101011001100000", '1'), -- i=3042
      ("0100011001100000", '-'), -- i=3043
      ("0000011010010101", '-'), -- i=3044
      ("1000011001100011", '-'), -- i=3045
      ("1001011001100011", '-'), -- i=3046
      ("1010011001100011", '-'), -- i=3047
      ("1011011001100011", '-'), -- i=3048
      ("0101011001100000", '1'), -- i=3049
      ("0100011001100000", '-'), -- i=3050
      ("0000011000100111", '-'), -- i=3051
      ("1000011001100100", '-'), -- i=3052
      ("1001011001100100", '-'), -- i=3053
      ("1010011001100100", '-'), -- i=3054
      ("1011011001100100", '-'), -- i=3055
      ("0101011001100000", '1'), -- i=3056
      ("0100011001100000", '-'), -- i=3057
      ("0000011000111010", '-'), -- i=3058
      ("1000011001100101", '-'), -- i=3059
      ("1001011001100101", '-'), -- i=3060
      ("1010011001100101", '-'), -- i=3061
      ("1011011001100101", '-'), -- i=3062
      ("0101011001100000", '1'), -- i=3063
      ("0100011001100000", '-'), -- i=3064
      ("0000011011101001", '-'), -- i=3065
      ("1000011001100110", '-'), -- i=3066
      ("1001011001100110", '-'), -- i=3067
      ("1010011001100110", '-'), -- i=3068
      ("1011011001100110", '-'), -- i=3069
      ("0101011001100000", '1'), -- i=3070
      ("0100011001100000", '-'), -- i=3071
      ("0000011010010101", '-'), -- i=3072
      ("1000011001100111", '-'), -- i=3073
      ("1001011001100111", '-'), -- i=3074
      ("1010011001100111", '-'), -- i=3075
      ("1011011001100111", '-'), -- i=3076
      ("0101011001100000", '1'), -- i=3077
      ("0100011001100000", '-'), -- i=3078
      ("0000011011011001", '-'), -- i=3079
      ("1000011001110000", '-'), -- i=3080
      ("1001011001110000", '-'), -- i=3081
      ("1010011001110000", '-'), -- i=3082
      ("1011011001110000", '-'), -- i=3083
      ("0101011001110000", '1'), -- i=3084
      ("0100011001110000", '-'), -- i=3085
      ("0000011001101111", '-'), -- i=3086
      ("1000011001110001", '-'), -- i=3087
      ("1001011001110001", '-'), -- i=3088
      ("1010011001110001", '-'), -- i=3089
      ("1011011001110001", '-'), -- i=3090
      ("0101011001110000", '1'), -- i=3091
      ("0100011001110000", '-'), -- i=3092
      ("0000011010011011", '-'), -- i=3093
      ("1000011001110010", '-'), -- i=3094
      ("1001011001110010", '-'), -- i=3095
      ("1010011001110010", '-'), -- i=3096
      ("1011011001110010", '-'), -- i=3097
      ("0101011001110000", '1'), -- i=3098
      ("0100011001110000", '-'), -- i=3099
      ("0000011011110101", '-'), -- i=3100
      ("1000011001110011", '-'), -- i=3101
      ("1001011001110011", '-'), -- i=3102
      ("1010011001110011", '-'), -- i=3103
      ("1011011001110011", '-'), -- i=3104
      ("0101011001110000", '1'), -- i=3105
      ("0100011001110000", '-'), -- i=3106
      ("0000011000000100", '-'), -- i=3107
      ("1000011001110100", '-'), -- i=3108
      ("1001011001110100", '-'), -- i=3109
      ("1010011001110100", '-'), -- i=3110
      ("1011011001110100", '-'), -- i=3111
      ("0101011001110000", '1'), -- i=3112
      ("0100011001110000", '-'), -- i=3113
      ("0000011001110111", '-'), -- i=3114
      ("1000011001110101", '-'), -- i=3115
      ("1001011001110101", '-'), -- i=3116
      ("1010011001110101", '-'), -- i=3117
      ("1011011001110101", '-'), -- i=3118
      ("0101011001110000", '1'), -- i=3119
      ("0100011001110000", '-'), -- i=3120
      ("0000011010000100", '-'), -- i=3121
      ("1000011001110110", '-'), -- i=3122
      ("1001011001110110", '-'), -- i=3123
      ("1010011001110110", '-'), -- i=3124
      ("1011011001110110", '-'), -- i=3125
      ("0101011001110000", '1'), -- i=3126
      ("0100011001110000", '-'), -- i=3127
      ("0000011000001001", '-'), -- i=3128
      ("1000011001110111", '-'), -- i=3129
      ("1001011001110111", '-'), -- i=3130
      ("1010011001110111", '-'), -- i=3131
      ("1011011001110111", '-'), -- i=3132
      ("0101011001110000", '1'), -- i=3133
      ("0100011001110000", '-'), -- i=3134
      ("0000011000001100", '-'), -- i=3135
      ("1000011100000000", '-'), -- i=3136
      ("1001011100000000", '-'), -- i=3137
      ("1010011100000000", '-'), -- i=3138
      ("1011011100000000", '-'), -- i=3139
      ("0101011100000000", '1'), -- i=3140
      ("0100011100000000", '-'), -- i=3141
      ("0000011110101101", '-'), -- i=3142
      ("1000011100000001", '-'), -- i=3143
      ("1001011100000001", '-'), -- i=3144
      ("1010011100000001", '-'), -- i=3145
      ("1011011100000001", '-'), -- i=3146
      ("0101011100000000", '1'), -- i=3147
      ("0100011100000000", '-'), -- i=3148
      ("0000011101000001", '-'), -- i=3149
      ("1000011100000010", '-'), -- i=3150
      ("1001011100000010", '-'), -- i=3151
      ("1010011100000010", '-'), -- i=3152
      ("1011011100000010", '-'), -- i=3153
      ("0101011100000000", '1'), -- i=3154
      ("0100011100000000", '-'), -- i=3155
      ("0000011110100010", '-'), -- i=3156
      ("1000011100000011", '-'), -- i=3157
      ("1001011100000011", '-'), -- i=3158
      ("1010011100000011", '-'), -- i=3159
      ("1011011100000011", '-'), -- i=3160
      ("0101011100000000", '1'), -- i=3161
      ("0100011100000000", '-'), -- i=3162
      ("0000011101011010", '-'), -- i=3163
      ("1000011100000100", '-'), -- i=3164
      ("1001011100000100", '-'), -- i=3165
      ("1010011100000100", '-'), -- i=3166
      ("1011011100000100", '-'), -- i=3167
      ("0101011100000000", '1'), -- i=3168
      ("0100011100000000", '-'), -- i=3169
      ("0000011111001100", '-'), -- i=3170
      ("1000011100000101", '-'), -- i=3171
      ("1001011100000101", '-'), -- i=3172
      ("1010011100000101", '-'), -- i=3173
      ("1011011100000101", '-'), -- i=3174
      ("0101011100000000", '1'), -- i=3175
      ("0100011100000000", '-'), -- i=3176
      ("0000011110000010", '-'), -- i=3177
      ("1000011100000110", '-'), -- i=3178
      ("1001011100000110", '-'), -- i=3179
      ("1010011100000110", '-'), -- i=3180
      ("1011011100000110", '-'), -- i=3181
      ("0101011100000000", '1'), -- i=3182
      ("0100011100000000", '-'), -- i=3183
      ("0000011111111010", '-'), -- i=3184
      ("1000011100000111", '-'), -- i=3185
      ("1001011100000111", '-'), -- i=3186
      ("1010011100000111", '-'), -- i=3187
      ("1011011100000111", '-'), -- i=3188
      ("0101011100000000", '1'), -- i=3189
      ("0100011100000000", '-'), -- i=3190
      ("0000011100001010", '-'), -- i=3191
      ("1000011100010000", '-'), -- i=3192
      ("1001011100010000", '-'), -- i=3193
      ("1010011100010000", '-'), -- i=3194
      ("1011011100010000", '-'), -- i=3195
      ("0101011100010000", '1'), -- i=3196
      ("0100011100010000", '-'), -- i=3197
      ("0000011111001000", '-'), -- i=3198
      ("1000011100010001", '-'), -- i=3199
      ("1001011100010001", '-'), -- i=3200
      ("1010011100010001", '-'), -- i=3201
      ("1011011100010001", '-'), -- i=3202
      ("0101011100010000", '1'), -- i=3203
      ("0100011100010000", '-'), -- i=3204
      ("0000011101111111", '-'), -- i=3205
      ("1000011100010010", '-'), -- i=3206
      ("1001011100010010", '-'), -- i=3207
      ("1010011100010010", '-'), -- i=3208
      ("1011011100010010", '-'), -- i=3209
      ("0101011100010000", '1'), -- i=3210
      ("0100011100010000", '-'), -- i=3211
      ("0000011101100101", '-'), -- i=3212
      ("1000011100010011", '-'), -- i=3213
      ("1001011100010011", '-'), -- i=3214
      ("1010011100010011", '-'), -- i=3215
      ("1011011100010011", '-'), -- i=3216
      ("0101011100010000", '1'), -- i=3217
      ("0100011100010000", '-'), -- i=3218
      ("0000011110001110", '-'), -- i=3219
      ("1000011100010100", '-'), -- i=3220
      ("1001011100010100", '-'), -- i=3221
      ("1010011100010100", '-'), -- i=3222
      ("1011011100010100", '-'), -- i=3223
      ("0101011100010000", '1'), -- i=3224
      ("0100011100010000", '-'), -- i=3225
      ("0000011100001001", '-'), -- i=3226
      ("1000011100010101", '-'), -- i=3227
      ("1001011100010101", '-'), -- i=3228
      ("1010011100010101", '-'), -- i=3229
      ("1011011100010101", '-'), -- i=3230
      ("0101011100010000", '1'), -- i=3231
      ("0100011100010000", '-'), -- i=3232
      ("0000011111110010", '-'), -- i=3233
      ("1000011100010110", '-'), -- i=3234
      ("1001011100010110", '-'), -- i=3235
      ("1010011100010110", '-'), -- i=3236
      ("1011011100010110", '-'), -- i=3237
      ("0101011100010000", '1'), -- i=3238
      ("0100011100010000", '-'), -- i=3239
      ("0000011101010101", '-'), -- i=3240
      ("1000011100010111", '-'), -- i=3241
      ("1001011100010111", '-'), -- i=3242
      ("1010011100010111", '-'), -- i=3243
      ("1011011100010111", '-'), -- i=3244
      ("0101011100010000", '1'), -- i=3245
      ("0100011100010000", '-'), -- i=3246
      ("0000011100010100", '-'), -- i=3247
      ("1000011100100000", '-'), -- i=3248
      ("1001011100100000", '-'), -- i=3249
      ("1010011100100000", '-'), -- i=3250
      ("1011011100100000", '-'), -- i=3251
      ("0101011100100000", '1'), -- i=3252
      ("0100011100100000", '-'), -- i=3253
      ("0000011110010011", '-'), -- i=3254
      ("1000011100100001", '-'), -- i=3255
      ("1001011100100001", '-'), -- i=3256
      ("1010011100100001", '-'), -- i=3257
      ("1011011100100001", '-'), -- i=3258
      ("0101011100100000", '1'), -- i=3259
      ("0100011100100000", '-'), -- i=3260
      ("0000011110100000", '-'), -- i=3261
      ("1000011100100010", '-'), -- i=3262
      ("1001011100100010", '-'), -- i=3263
      ("1010011100100010", '-'), -- i=3264
      ("1011011100100010", '-'), -- i=3265
      ("0101011100100000", '1'), -- i=3266
      ("0100011100100000", '-'), -- i=3267
      ("0000011110010000", '-'), -- i=3268
      ("1000011100100011", '-'), -- i=3269
      ("1001011100100011", '-'), -- i=3270
      ("1010011100100011", '-'), -- i=3271
      ("1011011100100011", '-'), -- i=3272
      ("0101011100100000", '1'), -- i=3273
      ("0100011100100000", '-'), -- i=3274
      ("0000011110100111", '-'), -- i=3275
      ("1000011100100100", '-'), -- i=3276
      ("1001011100100100", '-'), -- i=3277
      ("1010011100100100", '-'), -- i=3278
      ("1011011100100100", '-'), -- i=3279
      ("0101011100100000", '1'), -- i=3280
      ("0100011100100000", '-'), -- i=3281
      ("0000011110011110", '-'), -- i=3282
      ("1000011100100101", '-'), -- i=3283
      ("1001011100100101", '-'), -- i=3284
      ("1010011100100101", '-'), -- i=3285
      ("1011011100100101", '-'), -- i=3286
      ("0101011100100000", '1'), -- i=3287
      ("0100011100100000", '-'), -- i=3288
      ("0000011101011000", '-'), -- i=3289
      ("1000011100100110", '-'), -- i=3290
      ("1001011100100110", '-'), -- i=3291
      ("1010011100100110", '-'), -- i=3292
      ("1011011100100110", '-'), -- i=3293
      ("0101011100100000", '1'), -- i=3294
      ("0100011100100000", '-'), -- i=3295
      ("0000011111101111", '-'), -- i=3296
      ("1000011100100111", '-'), -- i=3297
      ("1001011100100111", '-'), -- i=3298
      ("1010011100100111", '-'), -- i=3299
      ("1011011100100111", '-'), -- i=3300
      ("0101011100100000", '1'), -- i=3301
      ("0100011100100000", '-'), -- i=3302
      ("0000011101010000", '-'), -- i=3303
      ("1000011100110000", '-'), -- i=3304
      ("1001011100110000", '-'), -- i=3305
      ("1010011100110000", '-'), -- i=3306
      ("1011011100110000", '-'), -- i=3307
      ("0101011100110000", '1'), -- i=3308
      ("0100011100110000", '-'), -- i=3309
      ("0000011101010001", '-'), -- i=3310
      ("1000011100110001", '-'), -- i=3311
      ("1001011100110001", '-'), -- i=3312
      ("1010011100110001", '-'), -- i=3313
      ("1011011100110001", '-'), -- i=3314
      ("0101011100110000", '1'), -- i=3315
      ("0100011100110000", '-'), -- i=3316
      ("0000011101011110", '-'), -- i=3317
      ("1000011100110010", '-'), -- i=3318
      ("1001011100110010", '-'), -- i=3319
      ("1010011100110010", '-'), -- i=3320
      ("1011011100110010", '-'), -- i=3321
      ("0101011100110000", '1'), -- i=3322
      ("0100011100110000", '-'), -- i=3323
      ("0000011110000001", '-'), -- i=3324
      ("1000011100110011", '-'), -- i=3325
      ("1001011100110011", '-'), -- i=3326
      ("1010011100110011", '-'), -- i=3327
      ("1011011100110011", '-'), -- i=3328
      ("0101011100110000", '1'), -- i=3329
      ("0100011100110000", '-'), -- i=3330
      ("0000011100011110", '-'), -- i=3331
      ("1000011100110100", '-'), -- i=3332
      ("1001011100110100", '-'), -- i=3333
      ("1010011100110100", '-'), -- i=3334
      ("1011011100110100", '-'), -- i=3335
      ("0101011100110000", '1'), -- i=3336
      ("0100011100110000", '-'), -- i=3337
      ("0000011101010101", '-'), -- i=3338
      ("1000011100110101", '-'), -- i=3339
      ("1001011100110101", '-'), -- i=3340
      ("1010011100110101", '-'), -- i=3341
      ("1011011100110101", '-'), -- i=3342
      ("0101011100110000", '1'), -- i=3343
      ("0100011100110000", '-'), -- i=3344
      ("0000011110110110", '-'), -- i=3345
      ("1000011100110110", '-'), -- i=3346
      ("1001011100110110", '-'), -- i=3347
      ("1010011100110110", '-'), -- i=3348
      ("1011011100110110", '-'), -- i=3349
      ("0101011100110000", '1'), -- i=3350
      ("0100011100110000", '-'), -- i=3351
      ("0000011101011110", '-'), -- i=3352
      ("1000011100110111", '-'), -- i=3353
      ("1001011100110111", '-'), -- i=3354
      ("1010011100110111", '-'), -- i=3355
      ("1011011100110111", '-'), -- i=3356
      ("0101011100110000", '1'), -- i=3357
      ("0100011100110000", '-'), -- i=3358
      ("0000011111111100", '-'), -- i=3359
      ("1000011101000000", '-'), -- i=3360
      ("1001011101000000", '-'), -- i=3361
      ("1010011101000000", '-'), -- i=3362
      ("1011011101000000", '-'), -- i=3363
      ("0101011101000000", '1'), -- i=3364
      ("0100011101000000", '-'), -- i=3365
      ("0000011100110111", '-'), -- i=3366
      ("1000011101000001", '-'), -- i=3367
      ("1001011101000001", '-'), -- i=3368
      ("1010011101000001", '-'), -- i=3369
      ("1011011101000001", '-'), -- i=3370
      ("0101011101000000", '1'), -- i=3371
      ("0100011101000000", '-'), -- i=3372
      ("0000011101100110", '-'), -- i=3373
      ("1000011101000010", '-'), -- i=3374
      ("1001011101000010", '-'), -- i=3375
      ("1010011101000010", '-'), -- i=3376
      ("1011011101000010", '-'), -- i=3377
      ("0101011101000000", '1'), -- i=3378
      ("0100011101000000", '-'), -- i=3379
      ("0000011100010001", '-'), -- i=3380
      ("1000011101000011", '-'), -- i=3381
      ("1001011101000011", '-'), -- i=3382
      ("1010011101000011", '-'), -- i=3383
      ("1011011101000011", '-'), -- i=3384
      ("0101011101000000", '1'), -- i=3385
      ("0100011101000000", '-'), -- i=3386
      ("0000011101010100", '-'), -- i=3387
      ("1000011101000100", '-'), -- i=3388
      ("1001011101000100", '-'), -- i=3389
      ("1010011101000100", '-'), -- i=3390
      ("1011011101000100", '-'), -- i=3391
      ("0101011101000000", '1'), -- i=3392
      ("0100011101000000", '-'), -- i=3393
      ("0000011110100101", '-'), -- i=3394
      ("1000011101000101", '-'), -- i=3395
      ("1001011101000101", '-'), -- i=3396
      ("1010011101000101", '-'), -- i=3397
      ("1011011101000101", '-'), -- i=3398
      ("0101011101000000", '1'), -- i=3399
      ("0100011101000000", '-'), -- i=3400
      ("0000011111000100", '-'), -- i=3401
      ("1000011101000110", '-'), -- i=3402
      ("1001011101000110", '-'), -- i=3403
      ("1010011101000110", '-'), -- i=3404
      ("1011011101000110", '-'), -- i=3405
      ("0101011101000000", '1'), -- i=3406
      ("0100011101000000", '-'), -- i=3407
      ("0000011100000110", '-'), -- i=3408
      ("1000011101000111", '-'), -- i=3409
      ("1001011101000111", '-'), -- i=3410
      ("1010011101000111", '-'), -- i=3411
      ("1011011101000111", '-'), -- i=3412
      ("0101011101000000", '1'), -- i=3413
      ("0100011101000000", '-'), -- i=3414
      ("0000011100001100", '-'), -- i=3415
      ("1000011101010000", '-'), -- i=3416
      ("1001011101010000", '-'), -- i=3417
      ("1010011101010000", '-'), -- i=3418
      ("1011011101010000", '-'), -- i=3419
      ("0101011101010000", '1'), -- i=3420
      ("0100011101010000", '-'), -- i=3421
      ("0000011111011110", '-'), -- i=3422
      ("1000011101010001", '-'), -- i=3423
      ("1001011101010001", '-'), -- i=3424
      ("1010011101010001", '-'), -- i=3425
      ("1011011101010001", '-'), -- i=3426
      ("0101011101010000", '1'), -- i=3427
      ("0100011101010000", '-'), -- i=3428
      ("0000011100011011", '-'), -- i=3429
      ("1000011101010010", '-'), -- i=3430
      ("1001011101010010", '-'), -- i=3431
      ("1010011101010010", '-'), -- i=3432
      ("1011011101010010", '-'), -- i=3433
      ("0101011101010000", '1'), -- i=3434
      ("0100011101010000", '-'), -- i=3435
      ("0000011100001100", '-'), -- i=3436
      ("1000011101010011", '-'), -- i=3437
      ("1001011101010011", '-'), -- i=3438
      ("1010011101010011", '-'), -- i=3439
      ("1011011101010011", '-'), -- i=3440
      ("0101011101010000", '1'), -- i=3441
      ("0100011101010000", '-'), -- i=3442
      ("0000011100110110", '-'), -- i=3443
      ("1000011101010100", '-'), -- i=3444
      ("1001011101010100", '-'), -- i=3445
      ("1010011101010100", '-'), -- i=3446
      ("1011011101010100", '-'), -- i=3447
      ("0101011101010000", '1'), -- i=3448
      ("0100011101010000", '-'), -- i=3449
      ("0000011111010111", '-'), -- i=3450
      ("1000011101010101", '-'), -- i=3451
      ("1001011101010101", '-'), -- i=3452
      ("1010011101010101", '-'), -- i=3453
      ("1011011101010101", '-'), -- i=3454
      ("0101011101010000", '1'), -- i=3455
      ("0100011101010000", '-'), -- i=3456
      ("0000011110001110", '-'), -- i=3457
      ("1000011101010110", '-'), -- i=3458
      ("1001011101010110", '-'), -- i=3459
      ("1010011101010110", '-'), -- i=3460
      ("1011011101010110", '-'), -- i=3461
      ("0101011101010000", '1'), -- i=3462
      ("0100011101010000", '-'), -- i=3463
      ("0000011110010110", '-'), -- i=3464
      ("1000011101010111", '-'), -- i=3465
      ("1001011101010111", '-'), -- i=3466
      ("1010011101010111", '-'), -- i=3467
      ("1011011101010111", '-'), -- i=3468
      ("0101011101010000", '1'), -- i=3469
      ("0100011101010000", '-'), -- i=3470
      ("0000011110111110", '-'), -- i=3471
      ("1000011101100000", '-'), -- i=3472
      ("1001011101100000", '-'), -- i=3473
      ("1010011101100000", '-'), -- i=3474
      ("1011011101100000", '-'), -- i=3475
      ("0101011101100000", '1'), -- i=3476
      ("0100011101100000", '-'), -- i=3477
      ("0000011111110011", '-'), -- i=3478
      ("1000011101100001", '-'), -- i=3479
      ("1001011101100001", '-'), -- i=3480
      ("1010011101100001", '-'), -- i=3481
      ("1011011101100001", '-'), -- i=3482
      ("0101011101100000", '1'), -- i=3483
      ("0100011101100000", '-'), -- i=3484
      ("0000011111010110", '-'), -- i=3485
      ("1000011101100010", '-'), -- i=3486
      ("1001011101100010", '-'), -- i=3487
      ("1010011101100010", '-'), -- i=3488
      ("1011011101100010", '-'), -- i=3489
      ("0101011101100000", '1'), -- i=3490
      ("0100011101100000", '-'), -- i=3491
      ("0000011100010111", '-'), -- i=3492
      ("1000011101100011", '-'), -- i=3493
      ("1001011101100011", '-'), -- i=3494
      ("1010011101100011", '-'), -- i=3495
      ("1011011101100011", '-'), -- i=3496
      ("0101011101100000", '1'), -- i=3497
      ("0100011101100000", '-'), -- i=3498
      ("0000011111001111", '-'), -- i=3499
      ("1000011101100100", '-'), -- i=3500
      ("1001011101100100", '-'), -- i=3501
      ("1010011101100100", '-'), -- i=3502
      ("1011011101100100", '-'), -- i=3503
      ("0101011101100000", '1'), -- i=3504
      ("0100011101100000", '-'), -- i=3505
      ("0000011101100010", '-'), -- i=3506
      ("1000011101100101", '-'), -- i=3507
      ("1001011101100101", '-'), -- i=3508
      ("1010011101100101", '-'), -- i=3509
      ("1011011101100101", '-'), -- i=3510
      ("0101011101100000", '1'), -- i=3511
      ("0100011101100000", '-'), -- i=3512
      ("0000011110110100", '-'), -- i=3513
      ("1000011101100110", '-'), -- i=3514
      ("1001011101100110", '-'), -- i=3515
      ("1010011101100110", '-'), -- i=3516
      ("1011011101100110", '-'), -- i=3517
      ("0101011101100000", '1'), -- i=3518
      ("0100011101100000", '-'), -- i=3519
      ("0000011101111100", '-'), -- i=3520
      ("1000011101100111", '-'), -- i=3521
      ("1001011101100111", '-'), -- i=3522
      ("1010011101100111", '-'), -- i=3523
      ("1011011101100111", '-'), -- i=3524
      ("0101011101100000", '1'), -- i=3525
      ("0100011101100000", '-'), -- i=3526
      ("0000011100110010", '-'), -- i=3527
      ("1000011101110000", '-'), -- i=3528
      ("1001011101110000", '-'), -- i=3529
      ("1010011101110000", '-'), -- i=3530
      ("1011011101110000", '-'), -- i=3531
      ("0101011101110000", '1'), -- i=3532
      ("0100011101110000", '-'), -- i=3533
      ("0000011110110000", '-'), -- i=3534
      ("1000011101110001", '-'), -- i=3535
      ("1001011101110001", '-'), -- i=3536
      ("1010011101110001", '-'), -- i=3537
      ("1011011101110001", '-'), -- i=3538
      ("0101011101110000", '1'), -- i=3539
      ("0100011101110000", '-'), -- i=3540
      ("0000011100011011", '-'), -- i=3541
      ("1000011101110010", '-'), -- i=3542
      ("1001011101110010", '-'), -- i=3543
      ("1010011101110010", '-'), -- i=3544
      ("1011011101110010", '-'), -- i=3545
      ("0101011101110000", '1'), -- i=3546
      ("0100011101110000", '-'), -- i=3547
      ("0000011110011100", '-'), -- i=3548
      ("1000011101110011", '-'), -- i=3549
      ("1001011101110011", '-'), -- i=3550
      ("1010011101110011", '-'), -- i=3551
      ("1011011101110011", '-'), -- i=3552
      ("0101011101110000", '1'), -- i=3553
      ("0100011101110000", '-'), -- i=3554
      ("0000011111011101", '-'), -- i=3555
      ("1000011101110100", '-'), -- i=3556
      ("1001011101110100", '-'), -- i=3557
      ("1010011101110100", '-'), -- i=3558
      ("1011011101110100", '-'), -- i=3559
      ("0101011101110000", '1'), -- i=3560
      ("0100011101110000", '-'), -- i=3561
      ("0000011100111110", '-'), -- i=3562
      ("1000011101110101", '-'), -- i=3563
      ("1001011101110101", '-'), -- i=3564
      ("1010011101110101", '-'), -- i=3565
      ("1011011101110101", '-'), -- i=3566
      ("0101011101110000", '1'), -- i=3567
      ("0100011101110000", '-'), -- i=3568
      ("0000011100000010", '-'), -- i=3569
      ("1000011101110110", '-'), -- i=3570
      ("1001011101110110", '-'), -- i=3571
      ("1010011101110110", '-'), -- i=3572
      ("1011011101110110", '-'), -- i=3573
      ("0101011101110000", '1'), -- i=3574
      ("0100011101110000", '-'), -- i=3575
      ("0000011100001000", '-'), -- i=3576
      ("1000011101110111", '-'), -- i=3577
      ("1001011101110111", '-'), -- i=3578
      ("1010011101110111", '-'), -- i=3579
      ("1011011101110111", '-'), -- i=3580
      ("0101011101110000", '1'), -- i=3581
      ("0100011101110000", '-'), -- i=3582
      ("0000011100001100", '-'));
  begin
    for i in patterns'range loop
      INST <= patterns(i).INST;
      wait for 10 ns;
      assert std_match(ALUOP, patterns(i).ALUOP) OR (ALUOP = "ZZ" AND patterns(i).ALUOP = "ZZ")
        report "wrong value for ALUOP, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).ALUOP) & ", found " & to_string(ALUOP) severity error;assert std_match(RS1, patterns(i).RS1) OR (RS1 = "ZZZ" AND patterns(i).RS1 = "ZZZ")
        report "wrong value for RS1, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).RS1) & ", found " & to_string(RS1) severity error;assert std_match(RS2, patterns(i).RS2) OR (RS2 = "ZZZ" AND patterns(i).RS2 = "ZZZ")
        report "wrong value for RS2, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).RS2) & ", found " & to_string(RS2) severity error;assert std_match(WS, patterns(i).WS) OR (WS = "ZZZ" AND patterns(i).WS = "ZZZ")
        report "wrong value for WS, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).WS) & ", found " & to_string(WS) severity error;assert std_match(STR, patterns(i).STR) OR (STR = 'Z' AND patterns(i).STR = 'Z')
        report "wrong value for STR, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).STR) & ", found " & std_logic'image(STR) severity error;assert std_match(WE, patterns(i).WE) OR (WE = 'Z' AND patterns(i).WE = 'Z')
        report "wrong value for WE, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).WE) & ", found " & std_logic'image(WE) severity error;assert std_match(DMUX, patterns(i).DMUX) OR (DMUX = "ZZ" AND patterns(i).DMUX = "ZZ")
        report "wrong value for DMUX, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).DMUX) & ", found " & to_string(DMUX) severity error;assert std_match(LDR, patterns(i).LDR) OR (LDR = 'Z' AND patterns(i).LDR = 'Z')
        report "wrong value for LDR, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).LDR) & ", found " & std_logic'image(LDR) severity error;end loop;
    wait;
  end process;
end behav;
