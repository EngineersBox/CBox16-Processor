--  A testbench for control_unit_RS2_tb
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity control_unit_RS2_tb is
end control_unit_RS2_tb;

architecture behav of control_unit_RS2_tb is
  component main
    port (
      INST: in std_logic_vector(15 downto 0);
      ALUOP: out std_logic_vector(1 downto 0);
      RS1: out std_logic_vector(2 downto 0);
      RS2: out std_logic_vector(2 downto 0);
      WS: out std_logic_vector(2 downto 0);
      STR: out std_logic;
      WE: out std_logic;
      DMUX: out std_logic_vector(1 downto 0);
      LDR: out std_logic);
  end component;

  signal INST : std_logic_vector(15 downto 0);
  signal ALUOP : std_logic_vector(1 downto 0);
  signal RS1 : std_logic_vector(2 downto 0);
  signal RS2 : std_logic_vector(2 downto 0);
  signal WS : std_logic_vector(2 downto 0);
  signal STR : std_logic;
  signal WE : std_logic;
  signal DMUX : std_logic_vector(1 downto 0);
  signal LDR : std_logic;
  function to_string ( a: std_logic_vector) return string is
      variable b : string (1 to a'length) := (others => NUL);
      variable stri : integer := 1; 
  begin
      for i in a'range loop
          b(stri) := std_logic'image(a((i)))(2);
      stri := stri+1;
      end loop;
      return b;
  end function;
begin
  main_0 : main port map (
    INST => INST,
    ALUOP => ALUOP,
    RS1 => RS1,
    RS2 => RS2,
    WS => WS,
    STR => STR,
    WE => WE,
    DMUX => DMUX,
    LDR => LDR );
  process
    type pattern_type is record
      INST : std_logic_vector(15 downto 0);
      RS2 : std_logic_vector(2 downto 0);
    end record;
    type pattern_array is array (natural range <>) of pattern_type;
    constant patterns : pattern_array := (
      ("1000000000000000", "000"), -- i=0
      ("1001000000000000", "000"), -- i=1
      ("1010000000000000", "000"), -- i=2
      ("1011000000000000", "000"), -- i=3
      ("0100000000000000", "000"), -- i=4
      ("1000000000000001", "001"), -- i=5
      ("1001000000000001", "001"), -- i=6
      ("1010000000000001", "001"), -- i=7
      ("1011000000000001", "001"), -- i=8
      ("0100000000000000", "000"), -- i=9
      ("1000000000000010", "010"), -- i=10
      ("1001000000000010", "010"), -- i=11
      ("1010000000000010", "010"), -- i=12
      ("1011000000000010", "010"), -- i=13
      ("0100000000000000", "000"), -- i=14
      ("1000000000000011", "011"), -- i=15
      ("1001000000000011", "011"), -- i=16
      ("1010000000000011", "011"), -- i=17
      ("1011000000000011", "011"), -- i=18
      ("0100000000000000", "000"), -- i=19
      ("1000000000000100", "100"), -- i=20
      ("1001000000000100", "100"), -- i=21
      ("1010000000000100", "100"), -- i=22
      ("1011000000000100", "100"), -- i=23
      ("0100000000000000", "000"), -- i=24
      ("1000000000000101", "101"), -- i=25
      ("1001000000000101", "101"), -- i=26
      ("1010000000000101", "101"), -- i=27
      ("1011000000000101", "101"), -- i=28
      ("0100000000000000", "000"), -- i=29
      ("1000000000000110", "110"), -- i=30
      ("1001000000000110", "110"), -- i=31
      ("1010000000000110", "110"), -- i=32
      ("1011000000000110", "110"), -- i=33
      ("0100000000000000", "000"), -- i=34
      ("1000000000000111", "111"), -- i=35
      ("1001000000000111", "111"), -- i=36
      ("1010000000000111", "111"), -- i=37
      ("1011000000000111", "111"), -- i=38
      ("0100000000000000", "000"), -- i=39
      ("1000000000010000", "000"), -- i=40
      ("1001000000010000", "000"), -- i=41
      ("1010000000010000", "000"), -- i=42
      ("1011000000010000", "000"), -- i=43
      ("0100000000010000", "000"), -- i=44
      ("1000000000010001", "001"), -- i=45
      ("1001000000010001", "001"), -- i=46
      ("1010000000010001", "001"), -- i=47
      ("1011000000010001", "001"), -- i=48
      ("0100000000010000", "000"), -- i=49
      ("1000000000010010", "010"), -- i=50
      ("1001000000010010", "010"), -- i=51
      ("1010000000010010", "010"), -- i=52
      ("1011000000010010", "010"), -- i=53
      ("0100000000010000", "000"), -- i=54
      ("1000000000010011", "011"), -- i=55
      ("1001000000010011", "011"), -- i=56
      ("1010000000010011", "011"), -- i=57
      ("1011000000010011", "011"), -- i=58
      ("0100000000010000", "000"), -- i=59
      ("1000000000010100", "100"), -- i=60
      ("1001000000010100", "100"), -- i=61
      ("1010000000010100", "100"), -- i=62
      ("1011000000010100", "100"), -- i=63
      ("0100000000010000", "000"), -- i=64
      ("1000000000010101", "101"), -- i=65
      ("1001000000010101", "101"), -- i=66
      ("1010000000010101", "101"), -- i=67
      ("1011000000010101", "101"), -- i=68
      ("0100000000010000", "000"), -- i=69
      ("1000000000010110", "110"), -- i=70
      ("1001000000010110", "110"), -- i=71
      ("1010000000010110", "110"), -- i=72
      ("1011000000010110", "110"), -- i=73
      ("0100000000010000", "000"), -- i=74
      ("1000000000010111", "111"), -- i=75
      ("1001000000010111", "111"), -- i=76
      ("1010000000010111", "111"), -- i=77
      ("1011000000010111", "111"), -- i=78
      ("0100000000010000", "000"), -- i=79
      ("1000000000100000", "000"), -- i=80
      ("1001000000100000", "000"), -- i=81
      ("1010000000100000", "000"), -- i=82
      ("1011000000100000", "000"), -- i=83
      ("0100000000100000", "000"), -- i=84
      ("1000000000100001", "001"), -- i=85
      ("1001000000100001", "001"), -- i=86
      ("1010000000100001", "001"), -- i=87
      ("1011000000100001", "001"), -- i=88
      ("0100000000100000", "000"), -- i=89
      ("1000000000100010", "010"), -- i=90
      ("1001000000100010", "010"), -- i=91
      ("1010000000100010", "010"), -- i=92
      ("1011000000100010", "010"), -- i=93
      ("0100000000100000", "000"), -- i=94
      ("1000000000100011", "011"), -- i=95
      ("1001000000100011", "011"), -- i=96
      ("1010000000100011", "011"), -- i=97
      ("1011000000100011", "011"), -- i=98
      ("0100000000100000", "000"), -- i=99
      ("1000000000100100", "100"), -- i=100
      ("1001000000100100", "100"), -- i=101
      ("1010000000100100", "100"), -- i=102
      ("1011000000100100", "100"), -- i=103
      ("0100000000100000", "000"), -- i=104
      ("1000000000100101", "101"), -- i=105
      ("1001000000100101", "101"), -- i=106
      ("1010000000100101", "101"), -- i=107
      ("1011000000100101", "101"), -- i=108
      ("0100000000100000", "000"), -- i=109
      ("1000000000100110", "110"), -- i=110
      ("1001000000100110", "110"), -- i=111
      ("1010000000100110", "110"), -- i=112
      ("1011000000100110", "110"), -- i=113
      ("0100000000100000", "000"), -- i=114
      ("1000000000100111", "111"), -- i=115
      ("1001000000100111", "111"), -- i=116
      ("1010000000100111", "111"), -- i=117
      ("1011000000100111", "111"), -- i=118
      ("0100000000100000", "000"), -- i=119
      ("1000000000110000", "000"), -- i=120
      ("1001000000110000", "000"), -- i=121
      ("1010000000110000", "000"), -- i=122
      ("1011000000110000", "000"), -- i=123
      ("0100000000110000", "000"), -- i=124
      ("1000000000110001", "001"), -- i=125
      ("1001000000110001", "001"), -- i=126
      ("1010000000110001", "001"), -- i=127
      ("1011000000110001", "001"), -- i=128
      ("0100000000110000", "000"), -- i=129
      ("1000000000110010", "010"), -- i=130
      ("1001000000110010", "010"), -- i=131
      ("1010000000110010", "010"), -- i=132
      ("1011000000110010", "010"), -- i=133
      ("0100000000110000", "000"), -- i=134
      ("1000000000110011", "011"), -- i=135
      ("1001000000110011", "011"), -- i=136
      ("1010000000110011", "011"), -- i=137
      ("1011000000110011", "011"), -- i=138
      ("0100000000110000", "000"), -- i=139
      ("1000000000110100", "100"), -- i=140
      ("1001000000110100", "100"), -- i=141
      ("1010000000110100", "100"), -- i=142
      ("1011000000110100", "100"), -- i=143
      ("0100000000110000", "000"), -- i=144
      ("1000000000110101", "101"), -- i=145
      ("1001000000110101", "101"), -- i=146
      ("1010000000110101", "101"), -- i=147
      ("1011000000110101", "101"), -- i=148
      ("0100000000110000", "000"), -- i=149
      ("1000000000110110", "110"), -- i=150
      ("1001000000110110", "110"), -- i=151
      ("1010000000110110", "110"), -- i=152
      ("1011000000110110", "110"), -- i=153
      ("0100000000110000", "000"), -- i=154
      ("1000000000110111", "111"), -- i=155
      ("1001000000110111", "111"), -- i=156
      ("1010000000110111", "111"), -- i=157
      ("1011000000110111", "111"), -- i=158
      ("0100000000110000", "000"), -- i=159
      ("1000000001000000", "000"), -- i=160
      ("1001000001000000", "000"), -- i=161
      ("1010000001000000", "000"), -- i=162
      ("1011000001000000", "000"), -- i=163
      ("0100000001000000", "000"), -- i=164
      ("1000000001000001", "001"), -- i=165
      ("1001000001000001", "001"), -- i=166
      ("1010000001000001", "001"), -- i=167
      ("1011000001000001", "001"), -- i=168
      ("0100000001000000", "000"), -- i=169
      ("1000000001000010", "010"), -- i=170
      ("1001000001000010", "010"), -- i=171
      ("1010000001000010", "010"), -- i=172
      ("1011000001000010", "010"), -- i=173
      ("0100000001000000", "000"), -- i=174
      ("1000000001000011", "011"), -- i=175
      ("1001000001000011", "011"), -- i=176
      ("1010000001000011", "011"), -- i=177
      ("1011000001000011", "011"), -- i=178
      ("0100000001000000", "000"), -- i=179
      ("1000000001000100", "100"), -- i=180
      ("1001000001000100", "100"), -- i=181
      ("1010000001000100", "100"), -- i=182
      ("1011000001000100", "100"), -- i=183
      ("0100000001000000", "000"), -- i=184
      ("1000000001000101", "101"), -- i=185
      ("1001000001000101", "101"), -- i=186
      ("1010000001000101", "101"), -- i=187
      ("1011000001000101", "101"), -- i=188
      ("0100000001000000", "000"), -- i=189
      ("1000000001000110", "110"), -- i=190
      ("1001000001000110", "110"), -- i=191
      ("1010000001000110", "110"), -- i=192
      ("1011000001000110", "110"), -- i=193
      ("0100000001000000", "000"), -- i=194
      ("1000000001000111", "111"), -- i=195
      ("1001000001000111", "111"), -- i=196
      ("1010000001000111", "111"), -- i=197
      ("1011000001000111", "111"), -- i=198
      ("0100000001000000", "000"), -- i=199
      ("1000000001010000", "000"), -- i=200
      ("1001000001010000", "000"), -- i=201
      ("1010000001010000", "000"), -- i=202
      ("1011000001010000", "000"), -- i=203
      ("0100000001010000", "000"), -- i=204
      ("1000000001010001", "001"), -- i=205
      ("1001000001010001", "001"), -- i=206
      ("1010000001010001", "001"), -- i=207
      ("1011000001010001", "001"), -- i=208
      ("0100000001010000", "000"), -- i=209
      ("1000000001010010", "010"), -- i=210
      ("1001000001010010", "010"), -- i=211
      ("1010000001010010", "010"), -- i=212
      ("1011000001010010", "010"), -- i=213
      ("0100000001010000", "000"), -- i=214
      ("1000000001010011", "011"), -- i=215
      ("1001000001010011", "011"), -- i=216
      ("1010000001010011", "011"), -- i=217
      ("1011000001010011", "011"), -- i=218
      ("0100000001010000", "000"), -- i=219
      ("1000000001010100", "100"), -- i=220
      ("1001000001010100", "100"), -- i=221
      ("1010000001010100", "100"), -- i=222
      ("1011000001010100", "100"), -- i=223
      ("0100000001010000", "000"), -- i=224
      ("1000000001010101", "101"), -- i=225
      ("1001000001010101", "101"), -- i=226
      ("1010000001010101", "101"), -- i=227
      ("1011000001010101", "101"), -- i=228
      ("0100000001010000", "000"), -- i=229
      ("1000000001010110", "110"), -- i=230
      ("1001000001010110", "110"), -- i=231
      ("1010000001010110", "110"), -- i=232
      ("1011000001010110", "110"), -- i=233
      ("0100000001010000", "000"), -- i=234
      ("1000000001010111", "111"), -- i=235
      ("1001000001010111", "111"), -- i=236
      ("1010000001010111", "111"), -- i=237
      ("1011000001010111", "111"), -- i=238
      ("0100000001010000", "000"), -- i=239
      ("1000000001100000", "000"), -- i=240
      ("1001000001100000", "000"), -- i=241
      ("1010000001100000", "000"), -- i=242
      ("1011000001100000", "000"), -- i=243
      ("0100000001100000", "000"), -- i=244
      ("1000000001100001", "001"), -- i=245
      ("1001000001100001", "001"), -- i=246
      ("1010000001100001", "001"), -- i=247
      ("1011000001100001", "001"), -- i=248
      ("0100000001100000", "000"), -- i=249
      ("1000000001100010", "010"), -- i=250
      ("1001000001100010", "010"), -- i=251
      ("1010000001100010", "010"), -- i=252
      ("1011000001100010", "010"), -- i=253
      ("0100000001100000", "000"), -- i=254
      ("1000000001100011", "011"), -- i=255
      ("1001000001100011", "011"), -- i=256
      ("1010000001100011", "011"), -- i=257
      ("1011000001100011", "011"), -- i=258
      ("0100000001100000", "000"), -- i=259
      ("1000000001100100", "100"), -- i=260
      ("1001000001100100", "100"), -- i=261
      ("1010000001100100", "100"), -- i=262
      ("1011000001100100", "100"), -- i=263
      ("0100000001100000", "000"), -- i=264
      ("1000000001100101", "101"), -- i=265
      ("1001000001100101", "101"), -- i=266
      ("1010000001100101", "101"), -- i=267
      ("1011000001100101", "101"), -- i=268
      ("0100000001100000", "000"), -- i=269
      ("1000000001100110", "110"), -- i=270
      ("1001000001100110", "110"), -- i=271
      ("1010000001100110", "110"), -- i=272
      ("1011000001100110", "110"), -- i=273
      ("0100000001100000", "000"), -- i=274
      ("1000000001100111", "111"), -- i=275
      ("1001000001100111", "111"), -- i=276
      ("1010000001100111", "111"), -- i=277
      ("1011000001100111", "111"), -- i=278
      ("0100000001100000", "000"), -- i=279
      ("1000000001110000", "000"), -- i=280
      ("1001000001110000", "000"), -- i=281
      ("1010000001110000", "000"), -- i=282
      ("1011000001110000", "000"), -- i=283
      ("0100000001110000", "000"), -- i=284
      ("1000000001110001", "001"), -- i=285
      ("1001000001110001", "001"), -- i=286
      ("1010000001110001", "001"), -- i=287
      ("1011000001110001", "001"), -- i=288
      ("0100000001110000", "000"), -- i=289
      ("1000000001110010", "010"), -- i=290
      ("1001000001110010", "010"), -- i=291
      ("1010000001110010", "010"), -- i=292
      ("1011000001110010", "010"), -- i=293
      ("0100000001110000", "000"), -- i=294
      ("1000000001110011", "011"), -- i=295
      ("1001000001110011", "011"), -- i=296
      ("1010000001110011", "011"), -- i=297
      ("1011000001110011", "011"), -- i=298
      ("0100000001110000", "000"), -- i=299
      ("1000000001110100", "100"), -- i=300
      ("1001000001110100", "100"), -- i=301
      ("1010000001110100", "100"), -- i=302
      ("1011000001110100", "100"), -- i=303
      ("0100000001110000", "000"), -- i=304
      ("1000000001110101", "101"), -- i=305
      ("1001000001110101", "101"), -- i=306
      ("1010000001110101", "101"), -- i=307
      ("1011000001110101", "101"), -- i=308
      ("0100000001110000", "000"), -- i=309
      ("1000000001110110", "110"), -- i=310
      ("1001000001110110", "110"), -- i=311
      ("1010000001110110", "110"), -- i=312
      ("1011000001110110", "110"), -- i=313
      ("0100000001110000", "000"), -- i=314
      ("1000000001110111", "111"), -- i=315
      ("1001000001110111", "111"), -- i=316
      ("1010000001110111", "111"), -- i=317
      ("1011000001110111", "111"), -- i=318
      ("0100000001110000", "000"), -- i=319
      ("1000000100000000", "000"), -- i=320
      ("1001000100000000", "000"), -- i=321
      ("1010000100000000", "000"), -- i=322
      ("1011000100000000", "000"), -- i=323
      ("0100000100000000", "001"), -- i=324
      ("1000000100000001", "001"), -- i=325
      ("1001000100000001", "001"), -- i=326
      ("1010000100000001", "001"), -- i=327
      ("1011000100000001", "001"), -- i=328
      ("0100000100000000", "001"), -- i=329
      ("1000000100000010", "010"), -- i=330
      ("1001000100000010", "010"), -- i=331
      ("1010000100000010", "010"), -- i=332
      ("1011000100000010", "010"), -- i=333
      ("0100000100000000", "001"), -- i=334
      ("1000000100000011", "011"), -- i=335
      ("1001000100000011", "011"), -- i=336
      ("1010000100000011", "011"), -- i=337
      ("1011000100000011", "011"), -- i=338
      ("0100000100000000", "001"), -- i=339
      ("1000000100000100", "100"), -- i=340
      ("1001000100000100", "100"), -- i=341
      ("1010000100000100", "100"), -- i=342
      ("1011000100000100", "100"), -- i=343
      ("0100000100000000", "001"), -- i=344
      ("1000000100000101", "101"), -- i=345
      ("1001000100000101", "101"), -- i=346
      ("1010000100000101", "101"), -- i=347
      ("1011000100000101", "101"), -- i=348
      ("0100000100000000", "001"), -- i=349
      ("1000000100000110", "110"), -- i=350
      ("1001000100000110", "110"), -- i=351
      ("1010000100000110", "110"), -- i=352
      ("1011000100000110", "110"), -- i=353
      ("0100000100000000", "001"), -- i=354
      ("1000000100000111", "111"), -- i=355
      ("1001000100000111", "111"), -- i=356
      ("1010000100000111", "111"), -- i=357
      ("1011000100000111", "111"), -- i=358
      ("0100000100000000", "001"), -- i=359
      ("1000000100010000", "000"), -- i=360
      ("1001000100010000", "000"), -- i=361
      ("1010000100010000", "000"), -- i=362
      ("1011000100010000", "000"), -- i=363
      ("0100000100010000", "001"), -- i=364
      ("1000000100010001", "001"), -- i=365
      ("1001000100010001", "001"), -- i=366
      ("1010000100010001", "001"), -- i=367
      ("1011000100010001", "001"), -- i=368
      ("0100000100010000", "001"), -- i=369
      ("1000000100010010", "010"), -- i=370
      ("1001000100010010", "010"), -- i=371
      ("1010000100010010", "010"), -- i=372
      ("1011000100010010", "010"), -- i=373
      ("0100000100010000", "001"), -- i=374
      ("1000000100010011", "011"), -- i=375
      ("1001000100010011", "011"), -- i=376
      ("1010000100010011", "011"), -- i=377
      ("1011000100010011", "011"), -- i=378
      ("0100000100010000", "001"), -- i=379
      ("1000000100010100", "100"), -- i=380
      ("1001000100010100", "100"), -- i=381
      ("1010000100010100", "100"), -- i=382
      ("1011000100010100", "100"), -- i=383
      ("0100000100010000", "001"), -- i=384
      ("1000000100010101", "101"), -- i=385
      ("1001000100010101", "101"), -- i=386
      ("1010000100010101", "101"), -- i=387
      ("1011000100010101", "101"), -- i=388
      ("0100000100010000", "001"), -- i=389
      ("1000000100010110", "110"), -- i=390
      ("1001000100010110", "110"), -- i=391
      ("1010000100010110", "110"), -- i=392
      ("1011000100010110", "110"), -- i=393
      ("0100000100010000", "001"), -- i=394
      ("1000000100010111", "111"), -- i=395
      ("1001000100010111", "111"), -- i=396
      ("1010000100010111", "111"), -- i=397
      ("1011000100010111", "111"), -- i=398
      ("0100000100010000", "001"), -- i=399
      ("1000000100100000", "000"), -- i=400
      ("1001000100100000", "000"), -- i=401
      ("1010000100100000", "000"), -- i=402
      ("1011000100100000", "000"), -- i=403
      ("0100000100100000", "001"), -- i=404
      ("1000000100100001", "001"), -- i=405
      ("1001000100100001", "001"), -- i=406
      ("1010000100100001", "001"), -- i=407
      ("1011000100100001", "001"), -- i=408
      ("0100000100100000", "001"), -- i=409
      ("1000000100100010", "010"), -- i=410
      ("1001000100100010", "010"), -- i=411
      ("1010000100100010", "010"), -- i=412
      ("1011000100100010", "010"), -- i=413
      ("0100000100100000", "001"), -- i=414
      ("1000000100100011", "011"), -- i=415
      ("1001000100100011", "011"), -- i=416
      ("1010000100100011", "011"), -- i=417
      ("1011000100100011", "011"), -- i=418
      ("0100000100100000", "001"), -- i=419
      ("1000000100100100", "100"), -- i=420
      ("1001000100100100", "100"), -- i=421
      ("1010000100100100", "100"), -- i=422
      ("1011000100100100", "100"), -- i=423
      ("0100000100100000", "001"), -- i=424
      ("1000000100100101", "101"), -- i=425
      ("1001000100100101", "101"), -- i=426
      ("1010000100100101", "101"), -- i=427
      ("1011000100100101", "101"), -- i=428
      ("0100000100100000", "001"), -- i=429
      ("1000000100100110", "110"), -- i=430
      ("1001000100100110", "110"), -- i=431
      ("1010000100100110", "110"), -- i=432
      ("1011000100100110", "110"), -- i=433
      ("0100000100100000", "001"), -- i=434
      ("1000000100100111", "111"), -- i=435
      ("1001000100100111", "111"), -- i=436
      ("1010000100100111", "111"), -- i=437
      ("1011000100100111", "111"), -- i=438
      ("0100000100100000", "001"), -- i=439
      ("1000000100110000", "000"), -- i=440
      ("1001000100110000", "000"), -- i=441
      ("1010000100110000", "000"), -- i=442
      ("1011000100110000", "000"), -- i=443
      ("0100000100110000", "001"), -- i=444
      ("1000000100110001", "001"), -- i=445
      ("1001000100110001", "001"), -- i=446
      ("1010000100110001", "001"), -- i=447
      ("1011000100110001", "001"), -- i=448
      ("0100000100110000", "001"), -- i=449
      ("1000000100110010", "010"), -- i=450
      ("1001000100110010", "010"), -- i=451
      ("1010000100110010", "010"), -- i=452
      ("1011000100110010", "010"), -- i=453
      ("0100000100110000", "001"), -- i=454
      ("1000000100110011", "011"), -- i=455
      ("1001000100110011", "011"), -- i=456
      ("1010000100110011", "011"), -- i=457
      ("1011000100110011", "011"), -- i=458
      ("0100000100110000", "001"), -- i=459
      ("1000000100110100", "100"), -- i=460
      ("1001000100110100", "100"), -- i=461
      ("1010000100110100", "100"), -- i=462
      ("1011000100110100", "100"), -- i=463
      ("0100000100110000", "001"), -- i=464
      ("1000000100110101", "101"), -- i=465
      ("1001000100110101", "101"), -- i=466
      ("1010000100110101", "101"), -- i=467
      ("1011000100110101", "101"), -- i=468
      ("0100000100110000", "001"), -- i=469
      ("1000000100110110", "110"), -- i=470
      ("1001000100110110", "110"), -- i=471
      ("1010000100110110", "110"), -- i=472
      ("1011000100110110", "110"), -- i=473
      ("0100000100110000", "001"), -- i=474
      ("1000000100110111", "111"), -- i=475
      ("1001000100110111", "111"), -- i=476
      ("1010000100110111", "111"), -- i=477
      ("1011000100110111", "111"), -- i=478
      ("0100000100110000", "001"), -- i=479
      ("1000000101000000", "000"), -- i=480
      ("1001000101000000", "000"), -- i=481
      ("1010000101000000", "000"), -- i=482
      ("1011000101000000", "000"), -- i=483
      ("0100000101000000", "001"), -- i=484
      ("1000000101000001", "001"), -- i=485
      ("1001000101000001", "001"), -- i=486
      ("1010000101000001", "001"), -- i=487
      ("1011000101000001", "001"), -- i=488
      ("0100000101000000", "001"), -- i=489
      ("1000000101000010", "010"), -- i=490
      ("1001000101000010", "010"), -- i=491
      ("1010000101000010", "010"), -- i=492
      ("1011000101000010", "010"), -- i=493
      ("0100000101000000", "001"), -- i=494
      ("1000000101000011", "011"), -- i=495
      ("1001000101000011", "011"), -- i=496
      ("1010000101000011", "011"), -- i=497
      ("1011000101000011", "011"), -- i=498
      ("0100000101000000", "001"), -- i=499
      ("1000000101000100", "100"), -- i=500
      ("1001000101000100", "100"), -- i=501
      ("1010000101000100", "100"), -- i=502
      ("1011000101000100", "100"), -- i=503
      ("0100000101000000", "001"), -- i=504
      ("1000000101000101", "101"), -- i=505
      ("1001000101000101", "101"), -- i=506
      ("1010000101000101", "101"), -- i=507
      ("1011000101000101", "101"), -- i=508
      ("0100000101000000", "001"), -- i=509
      ("1000000101000110", "110"), -- i=510
      ("1001000101000110", "110"), -- i=511
      ("1010000101000110", "110"), -- i=512
      ("1011000101000110", "110"), -- i=513
      ("0100000101000000", "001"), -- i=514
      ("1000000101000111", "111"), -- i=515
      ("1001000101000111", "111"), -- i=516
      ("1010000101000111", "111"), -- i=517
      ("1011000101000111", "111"), -- i=518
      ("0100000101000000", "001"), -- i=519
      ("1000000101010000", "000"), -- i=520
      ("1001000101010000", "000"), -- i=521
      ("1010000101010000", "000"), -- i=522
      ("1011000101010000", "000"), -- i=523
      ("0100000101010000", "001"), -- i=524
      ("1000000101010001", "001"), -- i=525
      ("1001000101010001", "001"), -- i=526
      ("1010000101010001", "001"), -- i=527
      ("1011000101010001", "001"), -- i=528
      ("0100000101010000", "001"), -- i=529
      ("1000000101010010", "010"), -- i=530
      ("1001000101010010", "010"), -- i=531
      ("1010000101010010", "010"), -- i=532
      ("1011000101010010", "010"), -- i=533
      ("0100000101010000", "001"), -- i=534
      ("1000000101010011", "011"), -- i=535
      ("1001000101010011", "011"), -- i=536
      ("1010000101010011", "011"), -- i=537
      ("1011000101010011", "011"), -- i=538
      ("0100000101010000", "001"), -- i=539
      ("1000000101010100", "100"), -- i=540
      ("1001000101010100", "100"), -- i=541
      ("1010000101010100", "100"), -- i=542
      ("1011000101010100", "100"), -- i=543
      ("0100000101010000", "001"), -- i=544
      ("1000000101010101", "101"), -- i=545
      ("1001000101010101", "101"), -- i=546
      ("1010000101010101", "101"), -- i=547
      ("1011000101010101", "101"), -- i=548
      ("0100000101010000", "001"), -- i=549
      ("1000000101010110", "110"), -- i=550
      ("1001000101010110", "110"), -- i=551
      ("1010000101010110", "110"), -- i=552
      ("1011000101010110", "110"), -- i=553
      ("0100000101010000", "001"), -- i=554
      ("1000000101010111", "111"), -- i=555
      ("1001000101010111", "111"), -- i=556
      ("1010000101010111", "111"), -- i=557
      ("1011000101010111", "111"), -- i=558
      ("0100000101010000", "001"), -- i=559
      ("1000000101100000", "000"), -- i=560
      ("1001000101100000", "000"), -- i=561
      ("1010000101100000", "000"), -- i=562
      ("1011000101100000", "000"), -- i=563
      ("0100000101100000", "001"), -- i=564
      ("1000000101100001", "001"), -- i=565
      ("1001000101100001", "001"), -- i=566
      ("1010000101100001", "001"), -- i=567
      ("1011000101100001", "001"), -- i=568
      ("0100000101100000", "001"), -- i=569
      ("1000000101100010", "010"), -- i=570
      ("1001000101100010", "010"), -- i=571
      ("1010000101100010", "010"), -- i=572
      ("1011000101100010", "010"), -- i=573
      ("0100000101100000", "001"), -- i=574
      ("1000000101100011", "011"), -- i=575
      ("1001000101100011", "011"), -- i=576
      ("1010000101100011", "011"), -- i=577
      ("1011000101100011", "011"), -- i=578
      ("0100000101100000", "001"), -- i=579
      ("1000000101100100", "100"), -- i=580
      ("1001000101100100", "100"), -- i=581
      ("1010000101100100", "100"), -- i=582
      ("1011000101100100", "100"), -- i=583
      ("0100000101100000", "001"), -- i=584
      ("1000000101100101", "101"), -- i=585
      ("1001000101100101", "101"), -- i=586
      ("1010000101100101", "101"), -- i=587
      ("1011000101100101", "101"), -- i=588
      ("0100000101100000", "001"), -- i=589
      ("1000000101100110", "110"), -- i=590
      ("1001000101100110", "110"), -- i=591
      ("1010000101100110", "110"), -- i=592
      ("1011000101100110", "110"), -- i=593
      ("0100000101100000", "001"), -- i=594
      ("1000000101100111", "111"), -- i=595
      ("1001000101100111", "111"), -- i=596
      ("1010000101100111", "111"), -- i=597
      ("1011000101100111", "111"), -- i=598
      ("0100000101100000", "001"), -- i=599
      ("1000000101110000", "000"), -- i=600
      ("1001000101110000", "000"), -- i=601
      ("1010000101110000", "000"), -- i=602
      ("1011000101110000", "000"), -- i=603
      ("0100000101110000", "001"), -- i=604
      ("1000000101110001", "001"), -- i=605
      ("1001000101110001", "001"), -- i=606
      ("1010000101110001", "001"), -- i=607
      ("1011000101110001", "001"), -- i=608
      ("0100000101110000", "001"), -- i=609
      ("1000000101110010", "010"), -- i=610
      ("1001000101110010", "010"), -- i=611
      ("1010000101110010", "010"), -- i=612
      ("1011000101110010", "010"), -- i=613
      ("0100000101110000", "001"), -- i=614
      ("1000000101110011", "011"), -- i=615
      ("1001000101110011", "011"), -- i=616
      ("1010000101110011", "011"), -- i=617
      ("1011000101110011", "011"), -- i=618
      ("0100000101110000", "001"), -- i=619
      ("1000000101110100", "100"), -- i=620
      ("1001000101110100", "100"), -- i=621
      ("1010000101110100", "100"), -- i=622
      ("1011000101110100", "100"), -- i=623
      ("0100000101110000", "001"), -- i=624
      ("1000000101110101", "101"), -- i=625
      ("1001000101110101", "101"), -- i=626
      ("1010000101110101", "101"), -- i=627
      ("1011000101110101", "101"), -- i=628
      ("0100000101110000", "001"), -- i=629
      ("1000000101110110", "110"), -- i=630
      ("1001000101110110", "110"), -- i=631
      ("1010000101110110", "110"), -- i=632
      ("1011000101110110", "110"), -- i=633
      ("0100000101110000", "001"), -- i=634
      ("1000000101110111", "111"), -- i=635
      ("1001000101110111", "111"), -- i=636
      ("1010000101110111", "111"), -- i=637
      ("1011000101110111", "111"), -- i=638
      ("0100000101110000", "001"), -- i=639
      ("1000001000000000", "000"), -- i=640
      ("1001001000000000", "000"), -- i=641
      ("1010001000000000", "000"), -- i=642
      ("1011001000000000", "000"), -- i=643
      ("0100001000000000", "010"), -- i=644
      ("1000001000000001", "001"), -- i=645
      ("1001001000000001", "001"), -- i=646
      ("1010001000000001", "001"), -- i=647
      ("1011001000000001", "001"), -- i=648
      ("0100001000000000", "010"), -- i=649
      ("1000001000000010", "010"), -- i=650
      ("1001001000000010", "010"), -- i=651
      ("1010001000000010", "010"), -- i=652
      ("1011001000000010", "010"), -- i=653
      ("0100001000000000", "010"), -- i=654
      ("1000001000000011", "011"), -- i=655
      ("1001001000000011", "011"), -- i=656
      ("1010001000000011", "011"), -- i=657
      ("1011001000000011", "011"), -- i=658
      ("0100001000000000", "010"), -- i=659
      ("1000001000000100", "100"), -- i=660
      ("1001001000000100", "100"), -- i=661
      ("1010001000000100", "100"), -- i=662
      ("1011001000000100", "100"), -- i=663
      ("0100001000000000", "010"), -- i=664
      ("1000001000000101", "101"), -- i=665
      ("1001001000000101", "101"), -- i=666
      ("1010001000000101", "101"), -- i=667
      ("1011001000000101", "101"), -- i=668
      ("0100001000000000", "010"), -- i=669
      ("1000001000000110", "110"), -- i=670
      ("1001001000000110", "110"), -- i=671
      ("1010001000000110", "110"), -- i=672
      ("1011001000000110", "110"), -- i=673
      ("0100001000000000", "010"), -- i=674
      ("1000001000000111", "111"), -- i=675
      ("1001001000000111", "111"), -- i=676
      ("1010001000000111", "111"), -- i=677
      ("1011001000000111", "111"), -- i=678
      ("0100001000000000", "010"), -- i=679
      ("1000001000010000", "000"), -- i=680
      ("1001001000010000", "000"), -- i=681
      ("1010001000010000", "000"), -- i=682
      ("1011001000010000", "000"), -- i=683
      ("0100001000010000", "010"), -- i=684
      ("1000001000010001", "001"), -- i=685
      ("1001001000010001", "001"), -- i=686
      ("1010001000010001", "001"), -- i=687
      ("1011001000010001", "001"), -- i=688
      ("0100001000010000", "010"), -- i=689
      ("1000001000010010", "010"), -- i=690
      ("1001001000010010", "010"), -- i=691
      ("1010001000010010", "010"), -- i=692
      ("1011001000010010", "010"), -- i=693
      ("0100001000010000", "010"), -- i=694
      ("1000001000010011", "011"), -- i=695
      ("1001001000010011", "011"), -- i=696
      ("1010001000010011", "011"), -- i=697
      ("1011001000010011", "011"), -- i=698
      ("0100001000010000", "010"), -- i=699
      ("1000001000010100", "100"), -- i=700
      ("1001001000010100", "100"), -- i=701
      ("1010001000010100", "100"), -- i=702
      ("1011001000010100", "100"), -- i=703
      ("0100001000010000", "010"), -- i=704
      ("1000001000010101", "101"), -- i=705
      ("1001001000010101", "101"), -- i=706
      ("1010001000010101", "101"), -- i=707
      ("1011001000010101", "101"), -- i=708
      ("0100001000010000", "010"), -- i=709
      ("1000001000010110", "110"), -- i=710
      ("1001001000010110", "110"), -- i=711
      ("1010001000010110", "110"), -- i=712
      ("1011001000010110", "110"), -- i=713
      ("0100001000010000", "010"), -- i=714
      ("1000001000010111", "111"), -- i=715
      ("1001001000010111", "111"), -- i=716
      ("1010001000010111", "111"), -- i=717
      ("1011001000010111", "111"), -- i=718
      ("0100001000010000", "010"), -- i=719
      ("1000001000100000", "000"), -- i=720
      ("1001001000100000", "000"), -- i=721
      ("1010001000100000", "000"), -- i=722
      ("1011001000100000", "000"), -- i=723
      ("0100001000100000", "010"), -- i=724
      ("1000001000100001", "001"), -- i=725
      ("1001001000100001", "001"), -- i=726
      ("1010001000100001", "001"), -- i=727
      ("1011001000100001", "001"), -- i=728
      ("0100001000100000", "010"), -- i=729
      ("1000001000100010", "010"), -- i=730
      ("1001001000100010", "010"), -- i=731
      ("1010001000100010", "010"), -- i=732
      ("1011001000100010", "010"), -- i=733
      ("0100001000100000", "010"), -- i=734
      ("1000001000100011", "011"), -- i=735
      ("1001001000100011", "011"), -- i=736
      ("1010001000100011", "011"), -- i=737
      ("1011001000100011", "011"), -- i=738
      ("0100001000100000", "010"), -- i=739
      ("1000001000100100", "100"), -- i=740
      ("1001001000100100", "100"), -- i=741
      ("1010001000100100", "100"), -- i=742
      ("1011001000100100", "100"), -- i=743
      ("0100001000100000", "010"), -- i=744
      ("1000001000100101", "101"), -- i=745
      ("1001001000100101", "101"), -- i=746
      ("1010001000100101", "101"), -- i=747
      ("1011001000100101", "101"), -- i=748
      ("0100001000100000", "010"), -- i=749
      ("1000001000100110", "110"), -- i=750
      ("1001001000100110", "110"), -- i=751
      ("1010001000100110", "110"), -- i=752
      ("1011001000100110", "110"), -- i=753
      ("0100001000100000", "010"), -- i=754
      ("1000001000100111", "111"), -- i=755
      ("1001001000100111", "111"), -- i=756
      ("1010001000100111", "111"), -- i=757
      ("1011001000100111", "111"), -- i=758
      ("0100001000100000", "010"), -- i=759
      ("1000001000110000", "000"), -- i=760
      ("1001001000110000", "000"), -- i=761
      ("1010001000110000", "000"), -- i=762
      ("1011001000110000", "000"), -- i=763
      ("0100001000110000", "010"), -- i=764
      ("1000001000110001", "001"), -- i=765
      ("1001001000110001", "001"), -- i=766
      ("1010001000110001", "001"), -- i=767
      ("1011001000110001", "001"), -- i=768
      ("0100001000110000", "010"), -- i=769
      ("1000001000110010", "010"), -- i=770
      ("1001001000110010", "010"), -- i=771
      ("1010001000110010", "010"), -- i=772
      ("1011001000110010", "010"), -- i=773
      ("0100001000110000", "010"), -- i=774
      ("1000001000110011", "011"), -- i=775
      ("1001001000110011", "011"), -- i=776
      ("1010001000110011", "011"), -- i=777
      ("1011001000110011", "011"), -- i=778
      ("0100001000110000", "010"), -- i=779
      ("1000001000110100", "100"), -- i=780
      ("1001001000110100", "100"), -- i=781
      ("1010001000110100", "100"), -- i=782
      ("1011001000110100", "100"), -- i=783
      ("0100001000110000", "010"), -- i=784
      ("1000001000110101", "101"), -- i=785
      ("1001001000110101", "101"), -- i=786
      ("1010001000110101", "101"), -- i=787
      ("1011001000110101", "101"), -- i=788
      ("0100001000110000", "010"), -- i=789
      ("1000001000110110", "110"), -- i=790
      ("1001001000110110", "110"), -- i=791
      ("1010001000110110", "110"), -- i=792
      ("1011001000110110", "110"), -- i=793
      ("0100001000110000", "010"), -- i=794
      ("1000001000110111", "111"), -- i=795
      ("1001001000110111", "111"), -- i=796
      ("1010001000110111", "111"), -- i=797
      ("1011001000110111", "111"), -- i=798
      ("0100001000110000", "010"), -- i=799
      ("1000001001000000", "000"), -- i=800
      ("1001001001000000", "000"), -- i=801
      ("1010001001000000", "000"), -- i=802
      ("1011001001000000", "000"), -- i=803
      ("0100001001000000", "010"), -- i=804
      ("1000001001000001", "001"), -- i=805
      ("1001001001000001", "001"), -- i=806
      ("1010001001000001", "001"), -- i=807
      ("1011001001000001", "001"), -- i=808
      ("0100001001000000", "010"), -- i=809
      ("1000001001000010", "010"), -- i=810
      ("1001001001000010", "010"), -- i=811
      ("1010001001000010", "010"), -- i=812
      ("1011001001000010", "010"), -- i=813
      ("0100001001000000", "010"), -- i=814
      ("1000001001000011", "011"), -- i=815
      ("1001001001000011", "011"), -- i=816
      ("1010001001000011", "011"), -- i=817
      ("1011001001000011", "011"), -- i=818
      ("0100001001000000", "010"), -- i=819
      ("1000001001000100", "100"), -- i=820
      ("1001001001000100", "100"), -- i=821
      ("1010001001000100", "100"), -- i=822
      ("1011001001000100", "100"), -- i=823
      ("0100001001000000", "010"), -- i=824
      ("1000001001000101", "101"), -- i=825
      ("1001001001000101", "101"), -- i=826
      ("1010001001000101", "101"), -- i=827
      ("1011001001000101", "101"), -- i=828
      ("0100001001000000", "010"), -- i=829
      ("1000001001000110", "110"), -- i=830
      ("1001001001000110", "110"), -- i=831
      ("1010001001000110", "110"), -- i=832
      ("1011001001000110", "110"), -- i=833
      ("0100001001000000", "010"), -- i=834
      ("1000001001000111", "111"), -- i=835
      ("1001001001000111", "111"), -- i=836
      ("1010001001000111", "111"), -- i=837
      ("1011001001000111", "111"), -- i=838
      ("0100001001000000", "010"), -- i=839
      ("1000001001010000", "000"), -- i=840
      ("1001001001010000", "000"), -- i=841
      ("1010001001010000", "000"), -- i=842
      ("1011001001010000", "000"), -- i=843
      ("0100001001010000", "010"), -- i=844
      ("1000001001010001", "001"), -- i=845
      ("1001001001010001", "001"), -- i=846
      ("1010001001010001", "001"), -- i=847
      ("1011001001010001", "001"), -- i=848
      ("0100001001010000", "010"), -- i=849
      ("1000001001010010", "010"), -- i=850
      ("1001001001010010", "010"), -- i=851
      ("1010001001010010", "010"), -- i=852
      ("1011001001010010", "010"), -- i=853
      ("0100001001010000", "010"), -- i=854
      ("1000001001010011", "011"), -- i=855
      ("1001001001010011", "011"), -- i=856
      ("1010001001010011", "011"), -- i=857
      ("1011001001010011", "011"), -- i=858
      ("0100001001010000", "010"), -- i=859
      ("1000001001010100", "100"), -- i=860
      ("1001001001010100", "100"), -- i=861
      ("1010001001010100", "100"), -- i=862
      ("1011001001010100", "100"), -- i=863
      ("0100001001010000", "010"), -- i=864
      ("1000001001010101", "101"), -- i=865
      ("1001001001010101", "101"), -- i=866
      ("1010001001010101", "101"), -- i=867
      ("1011001001010101", "101"), -- i=868
      ("0100001001010000", "010"), -- i=869
      ("1000001001010110", "110"), -- i=870
      ("1001001001010110", "110"), -- i=871
      ("1010001001010110", "110"), -- i=872
      ("1011001001010110", "110"), -- i=873
      ("0100001001010000", "010"), -- i=874
      ("1000001001010111", "111"), -- i=875
      ("1001001001010111", "111"), -- i=876
      ("1010001001010111", "111"), -- i=877
      ("1011001001010111", "111"), -- i=878
      ("0100001001010000", "010"), -- i=879
      ("1000001001100000", "000"), -- i=880
      ("1001001001100000", "000"), -- i=881
      ("1010001001100000", "000"), -- i=882
      ("1011001001100000", "000"), -- i=883
      ("0100001001100000", "010"), -- i=884
      ("1000001001100001", "001"), -- i=885
      ("1001001001100001", "001"), -- i=886
      ("1010001001100001", "001"), -- i=887
      ("1011001001100001", "001"), -- i=888
      ("0100001001100000", "010"), -- i=889
      ("1000001001100010", "010"), -- i=890
      ("1001001001100010", "010"), -- i=891
      ("1010001001100010", "010"), -- i=892
      ("1011001001100010", "010"), -- i=893
      ("0100001001100000", "010"), -- i=894
      ("1000001001100011", "011"), -- i=895
      ("1001001001100011", "011"), -- i=896
      ("1010001001100011", "011"), -- i=897
      ("1011001001100011", "011"), -- i=898
      ("0100001001100000", "010"), -- i=899
      ("1000001001100100", "100"), -- i=900
      ("1001001001100100", "100"), -- i=901
      ("1010001001100100", "100"), -- i=902
      ("1011001001100100", "100"), -- i=903
      ("0100001001100000", "010"), -- i=904
      ("1000001001100101", "101"), -- i=905
      ("1001001001100101", "101"), -- i=906
      ("1010001001100101", "101"), -- i=907
      ("1011001001100101", "101"), -- i=908
      ("0100001001100000", "010"), -- i=909
      ("1000001001100110", "110"), -- i=910
      ("1001001001100110", "110"), -- i=911
      ("1010001001100110", "110"), -- i=912
      ("1011001001100110", "110"), -- i=913
      ("0100001001100000", "010"), -- i=914
      ("1000001001100111", "111"), -- i=915
      ("1001001001100111", "111"), -- i=916
      ("1010001001100111", "111"), -- i=917
      ("1011001001100111", "111"), -- i=918
      ("0100001001100000", "010"), -- i=919
      ("1000001001110000", "000"), -- i=920
      ("1001001001110000", "000"), -- i=921
      ("1010001001110000", "000"), -- i=922
      ("1011001001110000", "000"), -- i=923
      ("0100001001110000", "010"), -- i=924
      ("1000001001110001", "001"), -- i=925
      ("1001001001110001", "001"), -- i=926
      ("1010001001110001", "001"), -- i=927
      ("1011001001110001", "001"), -- i=928
      ("0100001001110000", "010"), -- i=929
      ("1000001001110010", "010"), -- i=930
      ("1001001001110010", "010"), -- i=931
      ("1010001001110010", "010"), -- i=932
      ("1011001001110010", "010"), -- i=933
      ("0100001001110000", "010"), -- i=934
      ("1000001001110011", "011"), -- i=935
      ("1001001001110011", "011"), -- i=936
      ("1010001001110011", "011"), -- i=937
      ("1011001001110011", "011"), -- i=938
      ("0100001001110000", "010"), -- i=939
      ("1000001001110100", "100"), -- i=940
      ("1001001001110100", "100"), -- i=941
      ("1010001001110100", "100"), -- i=942
      ("1011001001110100", "100"), -- i=943
      ("0100001001110000", "010"), -- i=944
      ("1000001001110101", "101"), -- i=945
      ("1001001001110101", "101"), -- i=946
      ("1010001001110101", "101"), -- i=947
      ("1011001001110101", "101"), -- i=948
      ("0100001001110000", "010"), -- i=949
      ("1000001001110110", "110"), -- i=950
      ("1001001001110110", "110"), -- i=951
      ("1010001001110110", "110"), -- i=952
      ("1011001001110110", "110"), -- i=953
      ("0100001001110000", "010"), -- i=954
      ("1000001001110111", "111"), -- i=955
      ("1001001001110111", "111"), -- i=956
      ("1010001001110111", "111"), -- i=957
      ("1011001001110111", "111"), -- i=958
      ("0100001001110000", "010"), -- i=959
      ("1000001100000000", "000"), -- i=960
      ("1001001100000000", "000"), -- i=961
      ("1010001100000000", "000"), -- i=962
      ("1011001100000000", "000"), -- i=963
      ("0100001100000000", "011"), -- i=964
      ("1000001100000001", "001"), -- i=965
      ("1001001100000001", "001"), -- i=966
      ("1010001100000001", "001"), -- i=967
      ("1011001100000001", "001"), -- i=968
      ("0100001100000000", "011"), -- i=969
      ("1000001100000010", "010"), -- i=970
      ("1001001100000010", "010"), -- i=971
      ("1010001100000010", "010"), -- i=972
      ("1011001100000010", "010"), -- i=973
      ("0100001100000000", "011"), -- i=974
      ("1000001100000011", "011"), -- i=975
      ("1001001100000011", "011"), -- i=976
      ("1010001100000011", "011"), -- i=977
      ("1011001100000011", "011"), -- i=978
      ("0100001100000000", "011"), -- i=979
      ("1000001100000100", "100"), -- i=980
      ("1001001100000100", "100"), -- i=981
      ("1010001100000100", "100"), -- i=982
      ("1011001100000100", "100"), -- i=983
      ("0100001100000000", "011"), -- i=984
      ("1000001100000101", "101"), -- i=985
      ("1001001100000101", "101"), -- i=986
      ("1010001100000101", "101"), -- i=987
      ("1011001100000101", "101"), -- i=988
      ("0100001100000000", "011"), -- i=989
      ("1000001100000110", "110"), -- i=990
      ("1001001100000110", "110"), -- i=991
      ("1010001100000110", "110"), -- i=992
      ("1011001100000110", "110"), -- i=993
      ("0100001100000000", "011"), -- i=994
      ("1000001100000111", "111"), -- i=995
      ("1001001100000111", "111"), -- i=996
      ("1010001100000111", "111"), -- i=997
      ("1011001100000111", "111"), -- i=998
      ("0100001100000000", "011"), -- i=999
      ("1000001100010000", "000"), -- i=1000
      ("1001001100010000", "000"), -- i=1001
      ("1010001100010000", "000"), -- i=1002
      ("1011001100010000", "000"), -- i=1003
      ("0100001100010000", "011"), -- i=1004
      ("1000001100010001", "001"), -- i=1005
      ("1001001100010001", "001"), -- i=1006
      ("1010001100010001", "001"), -- i=1007
      ("1011001100010001", "001"), -- i=1008
      ("0100001100010000", "011"), -- i=1009
      ("1000001100010010", "010"), -- i=1010
      ("1001001100010010", "010"), -- i=1011
      ("1010001100010010", "010"), -- i=1012
      ("1011001100010010", "010"), -- i=1013
      ("0100001100010000", "011"), -- i=1014
      ("1000001100010011", "011"), -- i=1015
      ("1001001100010011", "011"), -- i=1016
      ("1010001100010011", "011"), -- i=1017
      ("1011001100010011", "011"), -- i=1018
      ("0100001100010000", "011"), -- i=1019
      ("1000001100010100", "100"), -- i=1020
      ("1001001100010100", "100"), -- i=1021
      ("1010001100010100", "100"), -- i=1022
      ("1011001100010100", "100"), -- i=1023
      ("0100001100010000", "011"), -- i=1024
      ("1000001100010101", "101"), -- i=1025
      ("1001001100010101", "101"), -- i=1026
      ("1010001100010101", "101"), -- i=1027
      ("1011001100010101", "101"), -- i=1028
      ("0100001100010000", "011"), -- i=1029
      ("1000001100010110", "110"), -- i=1030
      ("1001001100010110", "110"), -- i=1031
      ("1010001100010110", "110"), -- i=1032
      ("1011001100010110", "110"), -- i=1033
      ("0100001100010000", "011"), -- i=1034
      ("1000001100010111", "111"), -- i=1035
      ("1001001100010111", "111"), -- i=1036
      ("1010001100010111", "111"), -- i=1037
      ("1011001100010111", "111"), -- i=1038
      ("0100001100010000", "011"), -- i=1039
      ("1000001100100000", "000"), -- i=1040
      ("1001001100100000", "000"), -- i=1041
      ("1010001100100000", "000"), -- i=1042
      ("1011001100100000", "000"), -- i=1043
      ("0100001100100000", "011"), -- i=1044
      ("1000001100100001", "001"), -- i=1045
      ("1001001100100001", "001"), -- i=1046
      ("1010001100100001", "001"), -- i=1047
      ("1011001100100001", "001"), -- i=1048
      ("0100001100100000", "011"), -- i=1049
      ("1000001100100010", "010"), -- i=1050
      ("1001001100100010", "010"), -- i=1051
      ("1010001100100010", "010"), -- i=1052
      ("1011001100100010", "010"), -- i=1053
      ("0100001100100000", "011"), -- i=1054
      ("1000001100100011", "011"), -- i=1055
      ("1001001100100011", "011"), -- i=1056
      ("1010001100100011", "011"), -- i=1057
      ("1011001100100011", "011"), -- i=1058
      ("0100001100100000", "011"), -- i=1059
      ("1000001100100100", "100"), -- i=1060
      ("1001001100100100", "100"), -- i=1061
      ("1010001100100100", "100"), -- i=1062
      ("1011001100100100", "100"), -- i=1063
      ("0100001100100000", "011"), -- i=1064
      ("1000001100100101", "101"), -- i=1065
      ("1001001100100101", "101"), -- i=1066
      ("1010001100100101", "101"), -- i=1067
      ("1011001100100101", "101"), -- i=1068
      ("0100001100100000", "011"), -- i=1069
      ("1000001100100110", "110"), -- i=1070
      ("1001001100100110", "110"), -- i=1071
      ("1010001100100110", "110"), -- i=1072
      ("1011001100100110", "110"), -- i=1073
      ("0100001100100000", "011"), -- i=1074
      ("1000001100100111", "111"), -- i=1075
      ("1001001100100111", "111"), -- i=1076
      ("1010001100100111", "111"), -- i=1077
      ("1011001100100111", "111"), -- i=1078
      ("0100001100100000", "011"), -- i=1079
      ("1000001100110000", "000"), -- i=1080
      ("1001001100110000", "000"), -- i=1081
      ("1010001100110000", "000"), -- i=1082
      ("1011001100110000", "000"), -- i=1083
      ("0100001100110000", "011"), -- i=1084
      ("1000001100110001", "001"), -- i=1085
      ("1001001100110001", "001"), -- i=1086
      ("1010001100110001", "001"), -- i=1087
      ("1011001100110001", "001"), -- i=1088
      ("0100001100110000", "011"), -- i=1089
      ("1000001100110010", "010"), -- i=1090
      ("1001001100110010", "010"), -- i=1091
      ("1010001100110010", "010"), -- i=1092
      ("1011001100110010", "010"), -- i=1093
      ("0100001100110000", "011"), -- i=1094
      ("1000001100110011", "011"), -- i=1095
      ("1001001100110011", "011"), -- i=1096
      ("1010001100110011", "011"), -- i=1097
      ("1011001100110011", "011"), -- i=1098
      ("0100001100110000", "011"), -- i=1099
      ("1000001100110100", "100"), -- i=1100
      ("1001001100110100", "100"), -- i=1101
      ("1010001100110100", "100"), -- i=1102
      ("1011001100110100", "100"), -- i=1103
      ("0100001100110000", "011"), -- i=1104
      ("1000001100110101", "101"), -- i=1105
      ("1001001100110101", "101"), -- i=1106
      ("1010001100110101", "101"), -- i=1107
      ("1011001100110101", "101"), -- i=1108
      ("0100001100110000", "011"), -- i=1109
      ("1000001100110110", "110"), -- i=1110
      ("1001001100110110", "110"), -- i=1111
      ("1010001100110110", "110"), -- i=1112
      ("1011001100110110", "110"), -- i=1113
      ("0100001100110000", "011"), -- i=1114
      ("1000001100110111", "111"), -- i=1115
      ("1001001100110111", "111"), -- i=1116
      ("1010001100110111", "111"), -- i=1117
      ("1011001100110111", "111"), -- i=1118
      ("0100001100110000", "011"), -- i=1119
      ("1000001101000000", "000"), -- i=1120
      ("1001001101000000", "000"), -- i=1121
      ("1010001101000000", "000"), -- i=1122
      ("1011001101000000", "000"), -- i=1123
      ("0100001101000000", "011"), -- i=1124
      ("1000001101000001", "001"), -- i=1125
      ("1001001101000001", "001"), -- i=1126
      ("1010001101000001", "001"), -- i=1127
      ("1011001101000001", "001"), -- i=1128
      ("0100001101000000", "011"), -- i=1129
      ("1000001101000010", "010"), -- i=1130
      ("1001001101000010", "010"), -- i=1131
      ("1010001101000010", "010"), -- i=1132
      ("1011001101000010", "010"), -- i=1133
      ("0100001101000000", "011"), -- i=1134
      ("1000001101000011", "011"), -- i=1135
      ("1001001101000011", "011"), -- i=1136
      ("1010001101000011", "011"), -- i=1137
      ("1011001101000011", "011"), -- i=1138
      ("0100001101000000", "011"), -- i=1139
      ("1000001101000100", "100"), -- i=1140
      ("1001001101000100", "100"), -- i=1141
      ("1010001101000100", "100"), -- i=1142
      ("1011001101000100", "100"), -- i=1143
      ("0100001101000000", "011"), -- i=1144
      ("1000001101000101", "101"), -- i=1145
      ("1001001101000101", "101"), -- i=1146
      ("1010001101000101", "101"), -- i=1147
      ("1011001101000101", "101"), -- i=1148
      ("0100001101000000", "011"), -- i=1149
      ("1000001101000110", "110"), -- i=1150
      ("1001001101000110", "110"), -- i=1151
      ("1010001101000110", "110"), -- i=1152
      ("1011001101000110", "110"), -- i=1153
      ("0100001101000000", "011"), -- i=1154
      ("1000001101000111", "111"), -- i=1155
      ("1001001101000111", "111"), -- i=1156
      ("1010001101000111", "111"), -- i=1157
      ("1011001101000111", "111"), -- i=1158
      ("0100001101000000", "011"), -- i=1159
      ("1000001101010000", "000"), -- i=1160
      ("1001001101010000", "000"), -- i=1161
      ("1010001101010000", "000"), -- i=1162
      ("1011001101010000", "000"), -- i=1163
      ("0100001101010000", "011"), -- i=1164
      ("1000001101010001", "001"), -- i=1165
      ("1001001101010001", "001"), -- i=1166
      ("1010001101010001", "001"), -- i=1167
      ("1011001101010001", "001"), -- i=1168
      ("0100001101010000", "011"), -- i=1169
      ("1000001101010010", "010"), -- i=1170
      ("1001001101010010", "010"), -- i=1171
      ("1010001101010010", "010"), -- i=1172
      ("1011001101010010", "010"), -- i=1173
      ("0100001101010000", "011"), -- i=1174
      ("1000001101010011", "011"), -- i=1175
      ("1001001101010011", "011"), -- i=1176
      ("1010001101010011", "011"), -- i=1177
      ("1011001101010011", "011"), -- i=1178
      ("0100001101010000", "011"), -- i=1179
      ("1000001101010100", "100"), -- i=1180
      ("1001001101010100", "100"), -- i=1181
      ("1010001101010100", "100"), -- i=1182
      ("1011001101010100", "100"), -- i=1183
      ("0100001101010000", "011"), -- i=1184
      ("1000001101010101", "101"), -- i=1185
      ("1001001101010101", "101"), -- i=1186
      ("1010001101010101", "101"), -- i=1187
      ("1011001101010101", "101"), -- i=1188
      ("0100001101010000", "011"), -- i=1189
      ("1000001101010110", "110"), -- i=1190
      ("1001001101010110", "110"), -- i=1191
      ("1010001101010110", "110"), -- i=1192
      ("1011001101010110", "110"), -- i=1193
      ("0100001101010000", "011"), -- i=1194
      ("1000001101010111", "111"), -- i=1195
      ("1001001101010111", "111"), -- i=1196
      ("1010001101010111", "111"), -- i=1197
      ("1011001101010111", "111"), -- i=1198
      ("0100001101010000", "011"), -- i=1199
      ("1000001101100000", "000"), -- i=1200
      ("1001001101100000", "000"), -- i=1201
      ("1010001101100000", "000"), -- i=1202
      ("1011001101100000", "000"), -- i=1203
      ("0100001101100000", "011"), -- i=1204
      ("1000001101100001", "001"), -- i=1205
      ("1001001101100001", "001"), -- i=1206
      ("1010001101100001", "001"), -- i=1207
      ("1011001101100001", "001"), -- i=1208
      ("0100001101100000", "011"), -- i=1209
      ("1000001101100010", "010"), -- i=1210
      ("1001001101100010", "010"), -- i=1211
      ("1010001101100010", "010"), -- i=1212
      ("1011001101100010", "010"), -- i=1213
      ("0100001101100000", "011"), -- i=1214
      ("1000001101100011", "011"), -- i=1215
      ("1001001101100011", "011"), -- i=1216
      ("1010001101100011", "011"), -- i=1217
      ("1011001101100011", "011"), -- i=1218
      ("0100001101100000", "011"), -- i=1219
      ("1000001101100100", "100"), -- i=1220
      ("1001001101100100", "100"), -- i=1221
      ("1010001101100100", "100"), -- i=1222
      ("1011001101100100", "100"), -- i=1223
      ("0100001101100000", "011"), -- i=1224
      ("1000001101100101", "101"), -- i=1225
      ("1001001101100101", "101"), -- i=1226
      ("1010001101100101", "101"), -- i=1227
      ("1011001101100101", "101"), -- i=1228
      ("0100001101100000", "011"), -- i=1229
      ("1000001101100110", "110"), -- i=1230
      ("1001001101100110", "110"), -- i=1231
      ("1010001101100110", "110"), -- i=1232
      ("1011001101100110", "110"), -- i=1233
      ("0100001101100000", "011"), -- i=1234
      ("1000001101100111", "111"), -- i=1235
      ("1001001101100111", "111"), -- i=1236
      ("1010001101100111", "111"), -- i=1237
      ("1011001101100111", "111"), -- i=1238
      ("0100001101100000", "011"), -- i=1239
      ("1000001101110000", "000"), -- i=1240
      ("1001001101110000", "000"), -- i=1241
      ("1010001101110000", "000"), -- i=1242
      ("1011001101110000", "000"), -- i=1243
      ("0100001101110000", "011"), -- i=1244
      ("1000001101110001", "001"), -- i=1245
      ("1001001101110001", "001"), -- i=1246
      ("1010001101110001", "001"), -- i=1247
      ("1011001101110001", "001"), -- i=1248
      ("0100001101110000", "011"), -- i=1249
      ("1000001101110010", "010"), -- i=1250
      ("1001001101110010", "010"), -- i=1251
      ("1010001101110010", "010"), -- i=1252
      ("1011001101110010", "010"), -- i=1253
      ("0100001101110000", "011"), -- i=1254
      ("1000001101110011", "011"), -- i=1255
      ("1001001101110011", "011"), -- i=1256
      ("1010001101110011", "011"), -- i=1257
      ("1011001101110011", "011"), -- i=1258
      ("0100001101110000", "011"), -- i=1259
      ("1000001101110100", "100"), -- i=1260
      ("1001001101110100", "100"), -- i=1261
      ("1010001101110100", "100"), -- i=1262
      ("1011001101110100", "100"), -- i=1263
      ("0100001101110000", "011"), -- i=1264
      ("1000001101110101", "101"), -- i=1265
      ("1001001101110101", "101"), -- i=1266
      ("1010001101110101", "101"), -- i=1267
      ("1011001101110101", "101"), -- i=1268
      ("0100001101110000", "011"), -- i=1269
      ("1000001101110110", "110"), -- i=1270
      ("1001001101110110", "110"), -- i=1271
      ("1010001101110110", "110"), -- i=1272
      ("1011001101110110", "110"), -- i=1273
      ("0100001101110000", "011"), -- i=1274
      ("1000001101110111", "111"), -- i=1275
      ("1001001101110111", "111"), -- i=1276
      ("1010001101110111", "111"), -- i=1277
      ("1011001101110111", "111"), -- i=1278
      ("0100001101110000", "011"), -- i=1279
      ("1000010000000000", "000"), -- i=1280
      ("1001010000000000", "000"), -- i=1281
      ("1010010000000000", "000"), -- i=1282
      ("1011010000000000", "000"), -- i=1283
      ("0100010000000000", "100"), -- i=1284
      ("1000010000000001", "001"), -- i=1285
      ("1001010000000001", "001"), -- i=1286
      ("1010010000000001", "001"), -- i=1287
      ("1011010000000001", "001"), -- i=1288
      ("0100010000000000", "100"), -- i=1289
      ("1000010000000010", "010"), -- i=1290
      ("1001010000000010", "010"), -- i=1291
      ("1010010000000010", "010"), -- i=1292
      ("1011010000000010", "010"), -- i=1293
      ("0100010000000000", "100"), -- i=1294
      ("1000010000000011", "011"), -- i=1295
      ("1001010000000011", "011"), -- i=1296
      ("1010010000000011", "011"), -- i=1297
      ("1011010000000011", "011"), -- i=1298
      ("0100010000000000", "100"), -- i=1299
      ("1000010000000100", "100"), -- i=1300
      ("1001010000000100", "100"), -- i=1301
      ("1010010000000100", "100"), -- i=1302
      ("1011010000000100", "100"), -- i=1303
      ("0100010000000000", "100"), -- i=1304
      ("1000010000000101", "101"), -- i=1305
      ("1001010000000101", "101"), -- i=1306
      ("1010010000000101", "101"), -- i=1307
      ("1011010000000101", "101"), -- i=1308
      ("0100010000000000", "100"), -- i=1309
      ("1000010000000110", "110"), -- i=1310
      ("1001010000000110", "110"), -- i=1311
      ("1010010000000110", "110"), -- i=1312
      ("1011010000000110", "110"), -- i=1313
      ("0100010000000000", "100"), -- i=1314
      ("1000010000000111", "111"), -- i=1315
      ("1001010000000111", "111"), -- i=1316
      ("1010010000000111", "111"), -- i=1317
      ("1011010000000111", "111"), -- i=1318
      ("0100010000000000", "100"), -- i=1319
      ("1000010000010000", "000"), -- i=1320
      ("1001010000010000", "000"), -- i=1321
      ("1010010000010000", "000"), -- i=1322
      ("1011010000010000", "000"), -- i=1323
      ("0100010000010000", "100"), -- i=1324
      ("1000010000010001", "001"), -- i=1325
      ("1001010000010001", "001"), -- i=1326
      ("1010010000010001", "001"), -- i=1327
      ("1011010000010001", "001"), -- i=1328
      ("0100010000010000", "100"), -- i=1329
      ("1000010000010010", "010"), -- i=1330
      ("1001010000010010", "010"), -- i=1331
      ("1010010000010010", "010"), -- i=1332
      ("1011010000010010", "010"), -- i=1333
      ("0100010000010000", "100"), -- i=1334
      ("1000010000010011", "011"), -- i=1335
      ("1001010000010011", "011"), -- i=1336
      ("1010010000010011", "011"), -- i=1337
      ("1011010000010011", "011"), -- i=1338
      ("0100010000010000", "100"), -- i=1339
      ("1000010000010100", "100"), -- i=1340
      ("1001010000010100", "100"), -- i=1341
      ("1010010000010100", "100"), -- i=1342
      ("1011010000010100", "100"), -- i=1343
      ("0100010000010000", "100"), -- i=1344
      ("1000010000010101", "101"), -- i=1345
      ("1001010000010101", "101"), -- i=1346
      ("1010010000010101", "101"), -- i=1347
      ("1011010000010101", "101"), -- i=1348
      ("0100010000010000", "100"), -- i=1349
      ("1000010000010110", "110"), -- i=1350
      ("1001010000010110", "110"), -- i=1351
      ("1010010000010110", "110"), -- i=1352
      ("1011010000010110", "110"), -- i=1353
      ("0100010000010000", "100"), -- i=1354
      ("1000010000010111", "111"), -- i=1355
      ("1001010000010111", "111"), -- i=1356
      ("1010010000010111", "111"), -- i=1357
      ("1011010000010111", "111"), -- i=1358
      ("0100010000010000", "100"), -- i=1359
      ("1000010000100000", "000"), -- i=1360
      ("1001010000100000", "000"), -- i=1361
      ("1010010000100000", "000"), -- i=1362
      ("1011010000100000", "000"), -- i=1363
      ("0100010000100000", "100"), -- i=1364
      ("1000010000100001", "001"), -- i=1365
      ("1001010000100001", "001"), -- i=1366
      ("1010010000100001", "001"), -- i=1367
      ("1011010000100001", "001"), -- i=1368
      ("0100010000100000", "100"), -- i=1369
      ("1000010000100010", "010"), -- i=1370
      ("1001010000100010", "010"), -- i=1371
      ("1010010000100010", "010"), -- i=1372
      ("1011010000100010", "010"), -- i=1373
      ("0100010000100000", "100"), -- i=1374
      ("1000010000100011", "011"), -- i=1375
      ("1001010000100011", "011"), -- i=1376
      ("1010010000100011", "011"), -- i=1377
      ("1011010000100011", "011"), -- i=1378
      ("0100010000100000", "100"), -- i=1379
      ("1000010000100100", "100"), -- i=1380
      ("1001010000100100", "100"), -- i=1381
      ("1010010000100100", "100"), -- i=1382
      ("1011010000100100", "100"), -- i=1383
      ("0100010000100000", "100"), -- i=1384
      ("1000010000100101", "101"), -- i=1385
      ("1001010000100101", "101"), -- i=1386
      ("1010010000100101", "101"), -- i=1387
      ("1011010000100101", "101"), -- i=1388
      ("0100010000100000", "100"), -- i=1389
      ("1000010000100110", "110"), -- i=1390
      ("1001010000100110", "110"), -- i=1391
      ("1010010000100110", "110"), -- i=1392
      ("1011010000100110", "110"), -- i=1393
      ("0100010000100000", "100"), -- i=1394
      ("1000010000100111", "111"), -- i=1395
      ("1001010000100111", "111"), -- i=1396
      ("1010010000100111", "111"), -- i=1397
      ("1011010000100111", "111"), -- i=1398
      ("0100010000100000", "100"), -- i=1399
      ("1000010000110000", "000"), -- i=1400
      ("1001010000110000", "000"), -- i=1401
      ("1010010000110000", "000"), -- i=1402
      ("1011010000110000", "000"), -- i=1403
      ("0100010000110000", "100"), -- i=1404
      ("1000010000110001", "001"), -- i=1405
      ("1001010000110001", "001"), -- i=1406
      ("1010010000110001", "001"), -- i=1407
      ("1011010000110001", "001"), -- i=1408
      ("0100010000110000", "100"), -- i=1409
      ("1000010000110010", "010"), -- i=1410
      ("1001010000110010", "010"), -- i=1411
      ("1010010000110010", "010"), -- i=1412
      ("1011010000110010", "010"), -- i=1413
      ("0100010000110000", "100"), -- i=1414
      ("1000010000110011", "011"), -- i=1415
      ("1001010000110011", "011"), -- i=1416
      ("1010010000110011", "011"), -- i=1417
      ("1011010000110011", "011"), -- i=1418
      ("0100010000110000", "100"), -- i=1419
      ("1000010000110100", "100"), -- i=1420
      ("1001010000110100", "100"), -- i=1421
      ("1010010000110100", "100"), -- i=1422
      ("1011010000110100", "100"), -- i=1423
      ("0100010000110000", "100"), -- i=1424
      ("1000010000110101", "101"), -- i=1425
      ("1001010000110101", "101"), -- i=1426
      ("1010010000110101", "101"), -- i=1427
      ("1011010000110101", "101"), -- i=1428
      ("0100010000110000", "100"), -- i=1429
      ("1000010000110110", "110"), -- i=1430
      ("1001010000110110", "110"), -- i=1431
      ("1010010000110110", "110"), -- i=1432
      ("1011010000110110", "110"), -- i=1433
      ("0100010000110000", "100"), -- i=1434
      ("1000010000110111", "111"), -- i=1435
      ("1001010000110111", "111"), -- i=1436
      ("1010010000110111", "111"), -- i=1437
      ("1011010000110111", "111"), -- i=1438
      ("0100010000110000", "100"), -- i=1439
      ("1000010001000000", "000"), -- i=1440
      ("1001010001000000", "000"), -- i=1441
      ("1010010001000000", "000"), -- i=1442
      ("1011010001000000", "000"), -- i=1443
      ("0100010001000000", "100"), -- i=1444
      ("1000010001000001", "001"), -- i=1445
      ("1001010001000001", "001"), -- i=1446
      ("1010010001000001", "001"), -- i=1447
      ("1011010001000001", "001"), -- i=1448
      ("0100010001000000", "100"), -- i=1449
      ("1000010001000010", "010"), -- i=1450
      ("1001010001000010", "010"), -- i=1451
      ("1010010001000010", "010"), -- i=1452
      ("1011010001000010", "010"), -- i=1453
      ("0100010001000000", "100"), -- i=1454
      ("1000010001000011", "011"), -- i=1455
      ("1001010001000011", "011"), -- i=1456
      ("1010010001000011", "011"), -- i=1457
      ("1011010001000011", "011"), -- i=1458
      ("0100010001000000", "100"), -- i=1459
      ("1000010001000100", "100"), -- i=1460
      ("1001010001000100", "100"), -- i=1461
      ("1010010001000100", "100"), -- i=1462
      ("1011010001000100", "100"), -- i=1463
      ("0100010001000000", "100"), -- i=1464
      ("1000010001000101", "101"), -- i=1465
      ("1001010001000101", "101"), -- i=1466
      ("1010010001000101", "101"), -- i=1467
      ("1011010001000101", "101"), -- i=1468
      ("0100010001000000", "100"), -- i=1469
      ("1000010001000110", "110"), -- i=1470
      ("1001010001000110", "110"), -- i=1471
      ("1010010001000110", "110"), -- i=1472
      ("1011010001000110", "110"), -- i=1473
      ("0100010001000000", "100"), -- i=1474
      ("1000010001000111", "111"), -- i=1475
      ("1001010001000111", "111"), -- i=1476
      ("1010010001000111", "111"), -- i=1477
      ("1011010001000111", "111"), -- i=1478
      ("0100010001000000", "100"), -- i=1479
      ("1000010001010000", "000"), -- i=1480
      ("1001010001010000", "000"), -- i=1481
      ("1010010001010000", "000"), -- i=1482
      ("1011010001010000", "000"), -- i=1483
      ("0100010001010000", "100"), -- i=1484
      ("1000010001010001", "001"), -- i=1485
      ("1001010001010001", "001"), -- i=1486
      ("1010010001010001", "001"), -- i=1487
      ("1011010001010001", "001"), -- i=1488
      ("0100010001010000", "100"), -- i=1489
      ("1000010001010010", "010"), -- i=1490
      ("1001010001010010", "010"), -- i=1491
      ("1010010001010010", "010"), -- i=1492
      ("1011010001010010", "010"), -- i=1493
      ("0100010001010000", "100"), -- i=1494
      ("1000010001010011", "011"), -- i=1495
      ("1001010001010011", "011"), -- i=1496
      ("1010010001010011", "011"), -- i=1497
      ("1011010001010011", "011"), -- i=1498
      ("0100010001010000", "100"), -- i=1499
      ("1000010001010100", "100"), -- i=1500
      ("1001010001010100", "100"), -- i=1501
      ("1010010001010100", "100"), -- i=1502
      ("1011010001010100", "100"), -- i=1503
      ("0100010001010000", "100"), -- i=1504
      ("1000010001010101", "101"), -- i=1505
      ("1001010001010101", "101"), -- i=1506
      ("1010010001010101", "101"), -- i=1507
      ("1011010001010101", "101"), -- i=1508
      ("0100010001010000", "100"), -- i=1509
      ("1000010001010110", "110"), -- i=1510
      ("1001010001010110", "110"), -- i=1511
      ("1010010001010110", "110"), -- i=1512
      ("1011010001010110", "110"), -- i=1513
      ("0100010001010000", "100"), -- i=1514
      ("1000010001010111", "111"), -- i=1515
      ("1001010001010111", "111"), -- i=1516
      ("1010010001010111", "111"), -- i=1517
      ("1011010001010111", "111"), -- i=1518
      ("0100010001010000", "100"), -- i=1519
      ("1000010001100000", "000"), -- i=1520
      ("1001010001100000", "000"), -- i=1521
      ("1010010001100000", "000"), -- i=1522
      ("1011010001100000", "000"), -- i=1523
      ("0100010001100000", "100"), -- i=1524
      ("1000010001100001", "001"), -- i=1525
      ("1001010001100001", "001"), -- i=1526
      ("1010010001100001", "001"), -- i=1527
      ("1011010001100001", "001"), -- i=1528
      ("0100010001100000", "100"), -- i=1529
      ("1000010001100010", "010"), -- i=1530
      ("1001010001100010", "010"), -- i=1531
      ("1010010001100010", "010"), -- i=1532
      ("1011010001100010", "010"), -- i=1533
      ("0100010001100000", "100"), -- i=1534
      ("1000010001100011", "011"), -- i=1535
      ("1001010001100011", "011"), -- i=1536
      ("1010010001100011", "011"), -- i=1537
      ("1011010001100011", "011"), -- i=1538
      ("0100010001100000", "100"), -- i=1539
      ("1000010001100100", "100"), -- i=1540
      ("1001010001100100", "100"), -- i=1541
      ("1010010001100100", "100"), -- i=1542
      ("1011010001100100", "100"), -- i=1543
      ("0100010001100000", "100"), -- i=1544
      ("1000010001100101", "101"), -- i=1545
      ("1001010001100101", "101"), -- i=1546
      ("1010010001100101", "101"), -- i=1547
      ("1011010001100101", "101"), -- i=1548
      ("0100010001100000", "100"), -- i=1549
      ("1000010001100110", "110"), -- i=1550
      ("1001010001100110", "110"), -- i=1551
      ("1010010001100110", "110"), -- i=1552
      ("1011010001100110", "110"), -- i=1553
      ("0100010001100000", "100"), -- i=1554
      ("1000010001100111", "111"), -- i=1555
      ("1001010001100111", "111"), -- i=1556
      ("1010010001100111", "111"), -- i=1557
      ("1011010001100111", "111"), -- i=1558
      ("0100010001100000", "100"), -- i=1559
      ("1000010001110000", "000"), -- i=1560
      ("1001010001110000", "000"), -- i=1561
      ("1010010001110000", "000"), -- i=1562
      ("1011010001110000", "000"), -- i=1563
      ("0100010001110000", "100"), -- i=1564
      ("1000010001110001", "001"), -- i=1565
      ("1001010001110001", "001"), -- i=1566
      ("1010010001110001", "001"), -- i=1567
      ("1011010001110001", "001"), -- i=1568
      ("0100010001110000", "100"), -- i=1569
      ("1000010001110010", "010"), -- i=1570
      ("1001010001110010", "010"), -- i=1571
      ("1010010001110010", "010"), -- i=1572
      ("1011010001110010", "010"), -- i=1573
      ("0100010001110000", "100"), -- i=1574
      ("1000010001110011", "011"), -- i=1575
      ("1001010001110011", "011"), -- i=1576
      ("1010010001110011", "011"), -- i=1577
      ("1011010001110011", "011"), -- i=1578
      ("0100010001110000", "100"), -- i=1579
      ("1000010001110100", "100"), -- i=1580
      ("1001010001110100", "100"), -- i=1581
      ("1010010001110100", "100"), -- i=1582
      ("1011010001110100", "100"), -- i=1583
      ("0100010001110000", "100"), -- i=1584
      ("1000010001110101", "101"), -- i=1585
      ("1001010001110101", "101"), -- i=1586
      ("1010010001110101", "101"), -- i=1587
      ("1011010001110101", "101"), -- i=1588
      ("0100010001110000", "100"), -- i=1589
      ("1000010001110110", "110"), -- i=1590
      ("1001010001110110", "110"), -- i=1591
      ("1010010001110110", "110"), -- i=1592
      ("1011010001110110", "110"), -- i=1593
      ("0100010001110000", "100"), -- i=1594
      ("1000010001110111", "111"), -- i=1595
      ("1001010001110111", "111"), -- i=1596
      ("1010010001110111", "111"), -- i=1597
      ("1011010001110111", "111"), -- i=1598
      ("0100010001110000", "100"), -- i=1599
      ("1000010100000000", "000"), -- i=1600
      ("1001010100000000", "000"), -- i=1601
      ("1010010100000000", "000"), -- i=1602
      ("1011010100000000", "000"), -- i=1603
      ("0100010100000000", "101"), -- i=1604
      ("1000010100000001", "001"), -- i=1605
      ("1001010100000001", "001"), -- i=1606
      ("1010010100000001", "001"), -- i=1607
      ("1011010100000001", "001"), -- i=1608
      ("0100010100000000", "101"), -- i=1609
      ("1000010100000010", "010"), -- i=1610
      ("1001010100000010", "010"), -- i=1611
      ("1010010100000010", "010"), -- i=1612
      ("1011010100000010", "010"), -- i=1613
      ("0100010100000000", "101"), -- i=1614
      ("1000010100000011", "011"), -- i=1615
      ("1001010100000011", "011"), -- i=1616
      ("1010010100000011", "011"), -- i=1617
      ("1011010100000011", "011"), -- i=1618
      ("0100010100000000", "101"), -- i=1619
      ("1000010100000100", "100"), -- i=1620
      ("1001010100000100", "100"), -- i=1621
      ("1010010100000100", "100"), -- i=1622
      ("1011010100000100", "100"), -- i=1623
      ("0100010100000000", "101"), -- i=1624
      ("1000010100000101", "101"), -- i=1625
      ("1001010100000101", "101"), -- i=1626
      ("1010010100000101", "101"), -- i=1627
      ("1011010100000101", "101"), -- i=1628
      ("0100010100000000", "101"), -- i=1629
      ("1000010100000110", "110"), -- i=1630
      ("1001010100000110", "110"), -- i=1631
      ("1010010100000110", "110"), -- i=1632
      ("1011010100000110", "110"), -- i=1633
      ("0100010100000000", "101"), -- i=1634
      ("1000010100000111", "111"), -- i=1635
      ("1001010100000111", "111"), -- i=1636
      ("1010010100000111", "111"), -- i=1637
      ("1011010100000111", "111"), -- i=1638
      ("0100010100000000", "101"), -- i=1639
      ("1000010100010000", "000"), -- i=1640
      ("1001010100010000", "000"), -- i=1641
      ("1010010100010000", "000"), -- i=1642
      ("1011010100010000", "000"), -- i=1643
      ("0100010100010000", "101"), -- i=1644
      ("1000010100010001", "001"), -- i=1645
      ("1001010100010001", "001"), -- i=1646
      ("1010010100010001", "001"), -- i=1647
      ("1011010100010001", "001"), -- i=1648
      ("0100010100010000", "101"), -- i=1649
      ("1000010100010010", "010"), -- i=1650
      ("1001010100010010", "010"), -- i=1651
      ("1010010100010010", "010"), -- i=1652
      ("1011010100010010", "010"), -- i=1653
      ("0100010100010000", "101"), -- i=1654
      ("1000010100010011", "011"), -- i=1655
      ("1001010100010011", "011"), -- i=1656
      ("1010010100010011", "011"), -- i=1657
      ("1011010100010011", "011"), -- i=1658
      ("0100010100010000", "101"), -- i=1659
      ("1000010100010100", "100"), -- i=1660
      ("1001010100010100", "100"), -- i=1661
      ("1010010100010100", "100"), -- i=1662
      ("1011010100010100", "100"), -- i=1663
      ("0100010100010000", "101"), -- i=1664
      ("1000010100010101", "101"), -- i=1665
      ("1001010100010101", "101"), -- i=1666
      ("1010010100010101", "101"), -- i=1667
      ("1011010100010101", "101"), -- i=1668
      ("0100010100010000", "101"), -- i=1669
      ("1000010100010110", "110"), -- i=1670
      ("1001010100010110", "110"), -- i=1671
      ("1010010100010110", "110"), -- i=1672
      ("1011010100010110", "110"), -- i=1673
      ("0100010100010000", "101"), -- i=1674
      ("1000010100010111", "111"), -- i=1675
      ("1001010100010111", "111"), -- i=1676
      ("1010010100010111", "111"), -- i=1677
      ("1011010100010111", "111"), -- i=1678
      ("0100010100010000", "101"), -- i=1679
      ("1000010100100000", "000"), -- i=1680
      ("1001010100100000", "000"), -- i=1681
      ("1010010100100000", "000"), -- i=1682
      ("1011010100100000", "000"), -- i=1683
      ("0100010100100000", "101"), -- i=1684
      ("1000010100100001", "001"), -- i=1685
      ("1001010100100001", "001"), -- i=1686
      ("1010010100100001", "001"), -- i=1687
      ("1011010100100001", "001"), -- i=1688
      ("0100010100100000", "101"), -- i=1689
      ("1000010100100010", "010"), -- i=1690
      ("1001010100100010", "010"), -- i=1691
      ("1010010100100010", "010"), -- i=1692
      ("1011010100100010", "010"), -- i=1693
      ("0100010100100000", "101"), -- i=1694
      ("1000010100100011", "011"), -- i=1695
      ("1001010100100011", "011"), -- i=1696
      ("1010010100100011", "011"), -- i=1697
      ("1011010100100011", "011"), -- i=1698
      ("0100010100100000", "101"), -- i=1699
      ("1000010100100100", "100"), -- i=1700
      ("1001010100100100", "100"), -- i=1701
      ("1010010100100100", "100"), -- i=1702
      ("1011010100100100", "100"), -- i=1703
      ("0100010100100000", "101"), -- i=1704
      ("1000010100100101", "101"), -- i=1705
      ("1001010100100101", "101"), -- i=1706
      ("1010010100100101", "101"), -- i=1707
      ("1011010100100101", "101"), -- i=1708
      ("0100010100100000", "101"), -- i=1709
      ("1000010100100110", "110"), -- i=1710
      ("1001010100100110", "110"), -- i=1711
      ("1010010100100110", "110"), -- i=1712
      ("1011010100100110", "110"), -- i=1713
      ("0100010100100000", "101"), -- i=1714
      ("1000010100100111", "111"), -- i=1715
      ("1001010100100111", "111"), -- i=1716
      ("1010010100100111", "111"), -- i=1717
      ("1011010100100111", "111"), -- i=1718
      ("0100010100100000", "101"), -- i=1719
      ("1000010100110000", "000"), -- i=1720
      ("1001010100110000", "000"), -- i=1721
      ("1010010100110000", "000"), -- i=1722
      ("1011010100110000", "000"), -- i=1723
      ("0100010100110000", "101"), -- i=1724
      ("1000010100110001", "001"), -- i=1725
      ("1001010100110001", "001"), -- i=1726
      ("1010010100110001", "001"), -- i=1727
      ("1011010100110001", "001"), -- i=1728
      ("0100010100110000", "101"), -- i=1729
      ("1000010100110010", "010"), -- i=1730
      ("1001010100110010", "010"), -- i=1731
      ("1010010100110010", "010"), -- i=1732
      ("1011010100110010", "010"), -- i=1733
      ("0100010100110000", "101"), -- i=1734
      ("1000010100110011", "011"), -- i=1735
      ("1001010100110011", "011"), -- i=1736
      ("1010010100110011", "011"), -- i=1737
      ("1011010100110011", "011"), -- i=1738
      ("0100010100110000", "101"), -- i=1739
      ("1000010100110100", "100"), -- i=1740
      ("1001010100110100", "100"), -- i=1741
      ("1010010100110100", "100"), -- i=1742
      ("1011010100110100", "100"), -- i=1743
      ("0100010100110000", "101"), -- i=1744
      ("1000010100110101", "101"), -- i=1745
      ("1001010100110101", "101"), -- i=1746
      ("1010010100110101", "101"), -- i=1747
      ("1011010100110101", "101"), -- i=1748
      ("0100010100110000", "101"), -- i=1749
      ("1000010100110110", "110"), -- i=1750
      ("1001010100110110", "110"), -- i=1751
      ("1010010100110110", "110"), -- i=1752
      ("1011010100110110", "110"), -- i=1753
      ("0100010100110000", "101"), -- i=1754
      ("1000010100110111", "111"), -- i=1755
      ("1001010100110111", "111"), -- i=1756
      ("1010010100110111", "111"), -- i=1757
      ("1011010100110111", "111"), -- i=1758
      ("0100010100110000", "101"), -- i=1759
      ("1000010101000000", "000"), -- i=1760
      ("1001010101000000", "000"), -- i=1761
      ("1010010101000000", "000"), -- i=1762
      ("1011010101000000", "000"), -- i=1763
      ("0100010101000000", "101"), -- i=1764
      ("1000010101000001", "001"), -- i=1765
      ("1001010101000001", "001"), -- i=1766
      ("1010010101000001", "001"), -- i=1767
      ("1011010101000001", "001"), -- i=1768
      ("0100010101000000", "101"), -- i=1769
      ("1000010101000010", "010"), -- i=1770
      ("1001010101000010", "010"), -- i=1771
      ("1010010101000010", "010"), -- i=1772
      ("1011010101000010", "010"), -- i=1773
      ("0100010101000000", "101"), -- i=1774
      ("1000010101000011", "011"), -- i=1775
      ("1001010101000011", "011"), -- i=1776
      ("1010010101000011", "011"), -- i=1777
      ("1011010101000011", "011"), -- i=1778
      ("0100010101000000", "101"), -- i=1779
      ("1000010101000100", "100"), -- i=1780
      ("1001010101000100", "100"), -- i=1781
      ("1010010101000100", "100"), -- i=1782
      ("1011010101000100", "100"), -- i=1783
      ("0100010101000000", "101"), -- i=1784
      ("1000010101000101", "101"), -- i=1785
      ("1001010101000101", "101"), -- i=1786
      ("1010010101000101", "101"), -- i=1787
      ("1011010101000101", "101"), -- i=1788
      ("0100010101000000", "101"), -- i=1789
      ("1000010101000110", "110"), -- i=1790
      ("1001010101000110", "110"), -- i=1791
      ("1010010101000110", "110"), -- i=1792
      ("1011010101000110", "110"), -- i=1793
      ("0100010101000000", "101"), -- i=1794
      ("1000010101000111", "111"), -- i=1795
      ("1001010101000111", "111"), -- i=1796
      ("1010010101000111", "111"), -- i=1797
      ("1011010101000111", "111"), -- i=1798
      ("0100010101000000", "101"), -- i=1799
      ("1000010101010000", "000"), -- i=1800
      ("1001010101010000", "000"), -- i=1801
      ("1010010101010000", "000"), -- i=1802
      ("1011010101010000", "000"), -- i=1803
      ("0100010101010000", "101"), -- i=1804
      ("1000010101010001", "001"), -- i=1805
      ("1001010101010001", "001"), -- i=1806
      ("1010010101010001", "001"), -- i=1807
      ("1011010101010001", "001"), -- i=1808
      ("0100010101010000", "101"), -- i=1809
      ("1000010101010010", "010"), -- i=1810
      ("1001010101010010", "010"), -- i=1811
      ("1010010101010010", "010"), -- i=1812
      ("1011010101010010", "010"), -- i=1813
      ("0100010101010000", "101"), -- i=1814
      ("1000010101010011", "011"), -- i=1815
      ("1001010101010011", "011"), -- i=1816
      ("1010010101010011", "011"), -- i=1817
      ("1011010101010011", "011"), -- i=1818
      ("0100010101010000", "101"), -- i=1819
      ("1000010101010100", "100"), -- i=1820
      ("1001010101010100", "100"), -- i=1821
      ("1010010101010100", "100"), -- i=1822
      ("1011010101010100", "100"), -- i=1823
      ("0100010101010000", "101"), -- i=1824
      ("1000010101010101", "101"), -- i=1825
      ("1001010101010101", "101"), -- i=1826
      ("1010010101010101", "101"), -- i=1827
      ("1011010101010101", "101"), -- i=1828
      ("0100010101010000", "101"), -- i=1829
      ("1000010101010110", "110"), -- i=1830
      ("1001010101010110", "110"), -- i=1831
      ("1010010101010110", "110"), -- i=1832
      ("1011010101010110", "110"), -- i=1833
      ("0100010101010000", "101"), -- i=1834
      ("1000010101010111", "111"), -- i=1835
      ("1001010101010111", "111"), -- i=1836
      ("1010010101010111", "111"), -- i=1837
      ("1011010101010111", "111"), -- i=1838
      ("0100010101010000", "101"), -- i=1839
      ("1000010101100000", "000"), -- i=1840
      ("1001010101100000", "000"), -- i=1841
      ("1010010101100000", "000"), -- i=1842
      ("1011010101100000", "000"), -- i=1843
      ("0100010101100000", "101"), -- i=1844
      ("1000010101100001", "001"), -- i=1845
      ("1001010101100001", "001"), -- i=1846
      ("1010010101100001", "001"), -- i=1847
      ("1011010101100001", "001"), -- i=1848
      ("0100010101100000", "101"), -- i=1849
      ("1000010101100010", "010"), -- i=1850
      ("1001010101100010", "010"), -- i=1851
      ("1010010101100010", "010"), -- i=1852
      ("1011010101100010", "010"), -- i=1853
      ("0100010101100000", "101"), -- i=1854
      ("1000010101100011", "011"), -- i=1855
      ("1001010101100011", "011"), -- i=1856
      ("1010010101100011", "011"), -- i=1857
      ("1011010101100011", "011"), -- i=1858
      ("0100010101100000", "101"), -- i=1859
      ("1000010101100100", "100"), -- i=1860
      ("1001010101100100", "100"), -- i=1861
      ("1010010101100100", "100"), -- i=1862
      ("1011010101100100", "100"), -- i=1863
      ("0100010101100000", "101"), -- i=1864
      ("1000010101100101", "101"), -- i=1865
      ("1001010101100101", "101"), -- i=1866
      ("1010010101100101", "101"), -- i=1867
      ("1011010101100101", "101"), -- i=1868
      ("0100010101100000", "101"), -- i=1869
      ("1000010101100110", "110"), -- i=1870
      ("1001010101100110", "110"), -- i=1871
      ("1010010101100110", "110"), -- i=1872
      ("1011010101100110", "110"), -- i=1873
      ("0100010101100000", "101"), -- i=1874
      ("1000010101100111", "111"), -- i=1875
      ("1001010101100111", "111"), -- i=1876
      ("1010010101100111", "111"), -- i=1877
      ("1011010101100111", "111"), -- i=1878
      ("0100010101100000", "101"), -- i=1879
      ("1000010101110000", "000"), -- i=1880
      ("1001010101110000", "000"), -- i=1881
      ("1010010101110000", "000"), -- i=1882
      ("1011010101110000", "000"), -- i=1883
      ("0100010101110000", "101"), -- i=1884
      ("1000010101110001", "001"), -- i=1885
      ("1001010101110001", "001"), -- i=1886
      ("1010010101110001", "001"), -- i=1887
      ("1011010101110001", "001"), -- i=1888
      ("0100010101110000", "101"), -- i=1889
      ("1000010101110010", "010"), -- i=1890
      ("1001010101110010", "010"), -- i=1891
      ("1010010101110010", "010"), -- i=1892
      ("1011010101110010", "010"), -- i=1893
      ("0100010101110000", "101"), -- i=1894
      ("1000010101110011", "011"), -- i=1895
      ("1001010101110011", "011"), -- i=1896
      ("1010010101110011", "011"), -- i=1897
      ("1011010101110011", "011"), -- i=1898
      ("0100010101110000", "101"), -- i=1899
      ("1000010101110100", "100"), -- i=1900
      ("1001010101110100", "100"), -- i=1901
      ("1010010101110100", "100"), -- i=1902
      ("1011010101110100", "100"), -- i=1903
      ("0100010101110000", "101"), -- i=1904
      ("1000010101110101", "101"), -- i=1905
      ("1001010101110101", "101"), -- i=1906
      ("1010010101110101", "101"), -- i=1907
      ("1011010101110101", "101"), -- i=1908
      ("0100010101110000", "101"), -- i=1909
      ("1000010101110110", "110"), -- i=1910
      ("1001010101110110", "110"), -- i=1911
      ("1010010101110110", "110"), -- i=1912
      ("1011010101110110", "110"), -- i=1913
      ("0100010101110000", "101"), -- i=1914
      ("1000010101110111", "111"), -- i=1915
      ("1001010101110111", "111"), -- i=1916
      ("1010010101110111", "111"), -- i=1917
      ("1011010101110111", "111"), -- i=1918
      ("0100010101110000", "101"), -- i=1919
      ("1000011000000000", "000"), -- i=1920
      ("1001011000000000", "000"), -- i=1921
      ("1010011000000000", "000"), -- i=1922
      ("1011011000000000", "000"), -- i=1923
      ("0100011000000000", "110"), -- i=1924
      ("1000011000000001", "001"), -- i=1925
      ("1001011000000001", "001"), -- i=1926
      ("1010011000000001", "001"), -- i=1927
      ("1011011000000001", "001"), -- i=1928
      ("0100011000000000", "110"), -- i=1929
      ("1000011000000010", "010"), -- i=1930
      ("1001011000000010", "010"), -- i=1931
      ("1010011000000010", "010"), -- i=1932
      ("1011011000000010", "010"), -- i=1933
      ("0100011000000000", "110"), -- i=1934
      ("1000011000000011", "011"), -- i=1935
      ("1001011000000011", "011"), -- i=1936
      ("1010011000000011", "011"), -- i=1937
      ("1011011000000011", "011"), -- i=1938
      ("0100011000000000", "110"), -- i=1939
      ("1000011000000100", "100"), -- i=1940
      ("1001011000000100", "100"), -- i=1941
      ("1010011000000100", "100"), -- i=1942
      ("1011011000000100", "100"), -- i=1943
      ("0100011000000000", "110"), -- i=1944
      ("1000011000000101", "101"), -- i=1945
      ("1001011000000101", "101"), -- i=1946
      ("1010011000000101", "101"), -- i=1947
      ("1011011000000101", "101"), -- i=1948
      ("0100011000000000", "110"), -- i=1949
      ("1000011000000110", "110"), -- i=1950
      ("1001011000000110", "110"), -- i=1951
      ("1010011000000110", "110"), -- i=1952
      ("1011011000000110", "110"), -- i=1953
      ("0100011000000000", "110"), -- i=1954
      ("1000011000000111", "111"), -- i=1955
      ("1001011000000111", "111"), -- i=1956
      ("1010011000000111", "111"), -- i=1957
      ("1011011000000111", "111"), -- i=1958
      ("0100011000000000", "110"), -- i=1959
      ("1000011000010000", "000"), -- i=1960
      ("1001011000010000", "000"), -- i=1961
      ("1010011000010000", "000"), -- i=1962
      ("1011011000010000", "000"), -- i=1963
      ("0100011000010000", "110"), -- i=1964
      ("1000011000010001", "001"), -- i=1965
      ("1001011000010001", "001"), -- i=1966
      ("1010011000010001", "001"), -- i=1967
      ("1011011000010001", "001"), -- i=1968
      ("0100011000010000", "110"), -- i=1969
      ("1000011000010010", "010"), -- i=1970
      ("1001011000010010", "010"), -- i=1971
      ("1010011000010010", "010"), -- i=1972
      ("1011011000010010", "010"), -- i=1973
      ("0100011000010000", "110"), -- i=1974
      ("1000011000010011", "011"), -- i=1975
      ("1001011000010011", "011"), -- i=1976
      ("1010011000010011", "011"), -- i=1977
      ("1011011000010011", "011"), -- i=1978
      ("0100011000010000", "110"), -- i=1979
      ("1000011000010100", "100"), -- i=1980
      ("1001011000010100", "100"), -- i=1981
      ("1010011000010100", "100"), -- i=1982
      ("1011011000010100", "100"), -- i=1983
      ("0100011000010000", "110"), -- i=1984
      ("1000011000010101", "101"), -- i=1985
      ("1001011000010101", "101"), -- i=1986
      ("1010011000010101", "101"), -- i=1987
      ("1011011000010101", "101"), -- i=1988
      ("0100011000010000", "110"), -- i=1989
      ("1000011000010110", "110"), -- i=1990
      ("1001011000010110", "110"), -- i=1991
      ("1010011000010110", "110"), -- i=1992
      ("1011011000010110", "110"), -- i=1993
      ("0100011000010000", "110"), -- i=1994
      ("1000011000010111", "111"), -- i=1995
      ("1001011000010111", "111"), -- i=1996
      ("1010011000010111", "111"), -- i=1997
      ("1011011000010111", "111"), -- i=1998
      ("0100011000010000", "110"), -- i=1999
      ("1000011000100000", "000"), -- i=2000
      ("1001011000100000", "000"), -- i=2001
      ("1010011000100000", "000"), -- i=2002
      ("1011011000100000", "000"), -- i=2003
      ("0100011000100000", "110"), -- i=2004
      ("1000011000100001", "001"), -- i=2005
      ("1001011000100001", "001"), -- i=2006
      ("1010011000100001", "001"), -- i=2007
      ("1011011000100001", "001"), -- i=2008
      ("0100011000100000", "110"), -- i=2009
      ("1000011000100010", "010"), -- i=2010
      ("1001011000100010", "010"), -- i=2011
      ("1010011000100010", "010"), -- i=2012
      ("1011011000100010", "010"), -- i=2013
      ("0100011000100000", "110"), -- i=2014
      ("1000011000100011", "011"), -- i=2015
      ("1001011000100011", "011"), -- i=2016
      ("1010011000100011", "011"), -- i=2017
      ("1011011000100011", "011"), -- i=2018
      ("0100011000100000", "110"), -- i=2019
      ("1000011000100100", "100"), -- i=2020
      ("1001011000100100", "100"), -- i=2021
      ("1010011000100100", "100"), -- i=2022
      ("1011011000100100", "100"), -- i=2023
      ("0100011000100000", "110"), -- i=2024
      ("1000011000100101", "101"), -- i=2025
      ("1001011000100101", "101"), -- i=2026
      ("1010011000100101", "101"), -- i=2027
      ("1011011000100101", "101"), -- i=2028
      ("0100011000100000", "110"), -- i=2029
      ("1000011000100110", "110"), -- i=2030
      ("1001011000100110", "110"), -- i=2031
      ("1010011000100110", "110"), -- i=2032
      ("1011011000100110", "110"), -- i=2033
      ("0100011000100000", "110"), -- i=2034
      ("1000011000100111", "111"), -- i=2035
      ("1001011000100111", "111"), -- i=2036
      ("1010011000100111", "111"), -- i=2037
      ("1011011000100111", "111"), -- i=2038
      ("0100011000100000", "110"), -- i=2039
      ("1000011000110000", "000"), -- i=2040
      ("1001011000110000", "000"), -- i=2041
      ("1010011000110000", "000"), -- i=2042
      ("1011011000110000", "000"), -- i=2043
      ("0100011000110000", "110"), -- i=2044
      ("1000011000110001", "001"), -- i=2045
      ("1001011000110001", "001"), -- i=2046
      ("1010011000110001", "001"), -- i=2047
      ("1011011000110001", "001"), -- i=2048
      ("0100011000110000", "110"), -- i=2049
      ("1000011000110010", "010"), -- i=2050
      ("1001011000110010", "010"), -- i=2051
      ("1010011000110010", "010"), -- i=2052
      ("1011011000110010", "010"), -- i=2053
      ("0100011000110000", "110"), -- i=2054
      ("1000011000110011", "011"), -- i=2055
      ("1001011000110011", "011"), -- i=2056
      ("1010011000110011", "011"), -- i=2057
      ("1011011000110011", "011"), -- i=2058
      ("0100011000110000", "110"), -- i=2059
      ("1000011000110100", "100"), -- i=2060
      ("1001011000110100", "100"), -- i=2061
      ("1010011000110100", "100"), -- i=2062
      ("1011011000110100", "100"), -- i=2063
      ("0100011000110000", "110"), -- i=2064
      ("1000011000110101", "101"), -- i=2065
      ("1001011000110101", "101"), -- i=2066
      ("1010011000110101", "101"), -- i=2067
      ("1011011000110101", "101"), -- i=2068
      ("0100011000110000", "110"), -- i=2069
      ("1000011000110110", "110"), -- i=2070
      ("1001011000110110", "110"), -- i=2071
      ("1010011000110110", "110"), -- i=2072
      ("1011011000110110", "110"), -- i=2073
      ("0100011000110000", "110"), -- i=2074
      ("1000011000110111", "111"), -- i=2075
      ("1001011000110111", "111"), -- i=2076
      ("1010011000110111", "111"), -- i=2077
      ("1011011000110111", "111"), -- i=2078
      ("0100011000110000", "110"), -- i=2079
      ("1000011001000000", "000"), -- i=2080
      ("1001011001000000", "000"), -- i=2081
      ("1010011001000000", "000"), -- i=2082
      ("1011011001000000", "000"), -- i=2083
      ("0100011001000000", "110"), -- i=2084
      ("1000011001000001", "001"), -- i=2085
      ("1001011001000001", "001"), -- i=2086
      ("1010011001000001", "001"), -- i=2087
      ("1011011001000001", "001"), -- i=2088
      ("0100011001000000", "110"), -- i=2089
      ("1000011001000010", "010"), -- i=2090
      ("1001011001000010", "010"), -- i=2091
      ("1010011001000010", "010"), -- i=2092
      ("1011011001000010", "010"), -- i=2093
      ("0100011001000000", "110"), -- i=2094
      ("1000011001000011", "011"), -- i=2095
      ("1001011001000011", "011"), -- i=2096
      ("1010011001000011", "011"), -- i=2097
      ("1011011001000011", "011"), -- i=2098
      ("0100011001000000", "110"), -- i=2099
      ("1000011001000100", "100"), -- i=2100
      ("1001011001000100", "100"), -- i=2101
      ("1010011001000100", "100"), -- i=2102
      ("1011011001000100", "100"), -- i=2103
      ("0100011001000000", "110"), -- i=2104
      ("1000011001000101", "101"), -- i=2105
      ("1001011001000101", "101"), -- i=2106
      ("1010011001000101", "101"), -- i=2107
      ("1011011001000101", "101"), -- i=2108
      ("0100011001000000", "110"), -- i=2109
      ("1000011001000110", "110"), -- i=2110
      ("1001011001000110", "110"), -- i=2111
      ("1010011001000110", "110"), -- i=2112
      ("1011011001000110", "110"), -- i=2113
      ("0100011001000000", "110"), -- i=2114
      ("1000011001000111", "111"), -- i=2115
      ("1001011001000111", "111"), -- i=2116
      ("1010011001000111", "111"), -- i=2117
      ("1011011001000111", "111"), -- i=2118
      ("0100011001000000", "110"), -- i=2119
      ("1000011001010000", "000"), -- i=2120
      ("1001011001010000", "000"), -- i=2121
      ("1010011001010000", "000"), -- i=2122
      ("1011011001010000", "000"), -- i=2123
      ("0100011001010000", "110"), -- i=2124
      ("1000011001010001", "001"), -- i=2125
      ("1001011001010001", "001"), -- i=2126
      ("1010011001010001", "001"), -- i=2127
      ("1011011001010001", "001"), -- i=2128
      ("0100011001010000", "110"), -- i=2129
      ("1000011001010010", "010"), -- i=2130
      ("1001011001010010", "010"), -- i=2131
      ("1010011001010010", "010"), -- i=2132
      ("1011011001010010", "010"), -- i=2133
      ("0100011001010000", "110"), -- i=2134
      ("1000011001010011", "011"), -- i=2135
      ("1001011001010011", "011"), -- i=2136
      ("1010011001010011", "011"), -- i=2137
      ("1011011001010011", "011"), -- i=2138
      ("0100011001010000", "110"), -- i=2139
      ("1000011001010100", "100"), -- i=2140
      ("1001011001010100", "100"), -- i=2141
      ("1010011001010100", "100"), -- i=2142
      ("1011011001010100", "100"), -- i=2143
      ("0100011001010000", "110"), -- i=2144
      ("1000011001010101", "101"), -- i=2145
      ("1001011001010101", "101"), -- i=2146
      ("1010011001010101", "101"), -- i=2147
      ("1011011001010101", "101"), -- i=2148
      ("0100011001010000", "110"), -- i=2149
      ("1000011001010110", "110"), -- i=2150
      ("1001011001010110", "110"), -- i=2151
      ("1010011001010110", "110"), -- i=2152
      ("1011011001010110", "110"), -- i=2153
      ("0100011001010000", "110"), -- i=2154
      ("1000011001010111", "111"), -- i=2155
      ("1001011001010111", "111"), -- i=2156
      ("1010011001010111", "111"), -- i=2157
      ("1011011001010111", "111"), -- i=2158
      ("0100011001010000", "110"), -- i=2159
      ("1000011001100000", "000"), -- i=2160
      ("1001011001100000", "000"), -- i=2161
      ("1010011001100000", "000"), -- i=2162
      ("1011011001100000", "000"), -- i=2163
      ("0100011001100000", "110"), -- i=2164
      ("1000011001100001", "001"), -- i=2165
      ("1001011001100001", "001"), -- i=2166
      ("1010011001100001", "001"), -- i=2167
      ("1011011001100001", "001"), -- i=2168
      ("0100011001100000", "110"), -- i=2169
      ("1000011001100010", "010"), -- i=2170
      ("1001011001100010", "010"), -- i=2171
      ("1010011001100010", "010"), -- i=2172
      ("1011011001100010", "010"), -- i=2173
      ("0100011001100000", "110"), -- i=2174
      ("1000011001100011", "011"), -- i=2175
      ("1001011001100011", "011"), -- i=2176
      ("1010011001100011", "011"), -- i=2177
      ("1011011001100011", "011"), -- i=2178
      ("0100011001100000", "110"), -- i=2179
      ("1000011001100100", "100"), -- i=2180
      ("1001011001100100", "100"), -- i=2181
      ("1010011001100100", "100"), -- i=2182
      ("1011011001100100", "100"), -- i=2183
      ("0100011001100000", "110"), -- i=2184
      ("1000011001100101", "101"), -- i=2185
      ("1001011001100101", "101"), -- i=2186
      ("1010011001100101", "101"), -- i=2187
      ("1011011001100101", "101"), -- i=2188
      ("0100011001100000", "110"), -- i=2189
      ("1000011001100110", "110"), -- i=2190
      ("1001011001100110", "110"), -- i=2191
      ("1010011001100110", "110"), -- i=2192
      ("1011011001100110", "110"), -- i=2193
      ("0100011001100000", "110"), -- i=2194
      ("1000011001100111", "111"), -- i=2195
      ("1001011001100111", "111"), -- i=2196
      ("1010011001100111", "111"), -- i=2197
      ("1011011001100111", "111"), -- i=2198
      ("0100011001100000", "110"), -- i=2199
      ("1000011001110000", "000"), -- i=2200
      ("1001011001110000", "000"), -- i=2201
      ("1010011001110000", "000"), -- i=2202
      ("1011011001110000", "000"), -- i=2203
      ("0100011001110000", "110"), -- i=2204
      ("1000011001110001", "001"), -- i=2205
      ("1001011001110001", "001"), -- i=2206
      ("1010011001110001", "001"), -- i=2207
      ("1011011001110001", "001"), -- i=2208
      ("0100011001110000", "110"), -- i=2209
      ("1000011001110010", "010"), -- i=2210
      ("1001011001110010", "010"), -- i=2211
      ("1010011001110010", "010"), -- i=2212
      ("1011011001110010", "010"), -- i=2213
      ("0100011001110000", "110"), -- i=2214
      ("1000011001110011", "011"), -- i=2215
      ("1001011001110011", "011"), -- i=2216
      ("1010011001110011", "011"), -- i=2217
      ("1011011001110011", "011"), -- i=2218
      ("0100011001110000", "110"), -- i=2219
      ("1000011001110100", "100"), -- i=2220
      ("1001011001110100", "100"), -- i=2221
      ("1010011001110100", "100"), -- i=2222
      ("1011011001110100", "100"), -- i=2223
      ("0100011001110000", "110"), -- i=2224
      ("1000011001110101", "101"), -- i=2225
      ("1001011001110101", "101"), -- i=2226
      ("1010011001110101", "101"), -- i=2227
      ("1011011001110101", "101"), -- i=2228
      ("0100011001110000", "110"), -- i=2229
      ("1000011001110110", "110"), -- i=2230
      ("1001011001110110", "110"), -- i=2231
      ("1010011001110110", "110"), -- i=2232
      ("1011011001110110", "110"), -- i=2233
      ("0100011001110000", "110"), -- i=2234
      ("1000011001110111", "111"), -- i=2235
      ("1001011001110111", "111"), -- i=2236
      ("1010011001110111", "111"), -- i=2237
      ("1011011001110111", "111"), -- i=2238
      ("0100011001110000", "110"), -- i=2239
      ("1000011100000000", "000"), -- i=2240
      ("1001011100000000", "000"), -- i=2241
      ("1010011100000000", "000"), -- i=2242
      ("1011011100000000", "000"), -- i=2243
      ("0100011100000000", "111"), -- i=2244
      ("1000011100000001", "001"), -- i=2245
      ("1001011100000001", "001"), -- i=2246
      ("1010011100000001", "001"), -- i=2247
      ("1011011100000001", "001"), -- i=2248
      ("0100011100000000", "111"), -- i=2249
      ("1000011100000010", "010"), -- i=2250
      ("1001011100000010", "010"), -- i=2251
      ("1010011100000010", "010"), -- i=2252
      ("1011011100000010", "010"), -- i=2253
      ("0100011100000000", "111"), -- i=2254
      ("1000011100000011", "011"), -- i=2255
      ("1001011100000011", "011"), -- i=2256
      ("1010011100000011", "011"), -- i=2257
      ("1011011100000011", "011"), -- i=2258
      ("0100011100000000", "111"), -- i=2259
      ("1000011100000100", "100"), -- i=2260
      ("1001011100000100", "100"), -- i=2261
      ("1010011100000100", "100"), -- i=2262
      ("1011011100000100", "100"), -- i=2263
      ("0100011100000000", "111"), -- i=2264
      ("1000011100000101", "101"), -- i=2265
      ("1001011100000101", "101"), -- i=2266
      ("1010011100000101", "101"), -- i=2267
      ("1011011100000101", "101"), -- i=2268
      ("0100011100000000", "111"), -- i=2269
      ("1000011100000110", "110"), -- i=2270
      ("1001011100000110", "110"), -- i=2271
      ("1010011100000110", "110"), -- i=2272
      ("1011011100000110", "110"), -- i=2273
      ("0100011100000000", "111"), -- i=2274
      ("1000011100000111", "111"), -- i=2275
      ("1001011100000111", "111"), -- i=2276
      ("1010011100000111", "111"), -- i=2277
      ("1011011100000111", "111"), -- i=2278
      ("0100011100000000", "111"), -- i=2279
      ("1000011100010000", "000"), -- i=2280
      ("1001011100010000", "000"), -- i=2281
      ("1010011100010000", "000"), -- i=2282
      ("1011011100010000", "000"), -- i=2283
      ("0100011100010000", "111"), -- i=2284
      ("1000011100010001", "001"), -- i=2285
      ("1001011100010001", "001"), -- i=2286
      ("1010011100010001", "001"), -- i=2287
      ("1011011100010001", "001"), -- i=2288
      ("0100011100010000", "111"), -- i=2289
      ("1000011100010010", "010"), -- i=2290
      ("1001011100010010", "010"), -- i=2291
      ("1010011100010010", "010"), -- i=2292
      ("1011011100010010", "010"), -- i=2293
      ("0100011100010000", "111"), -- i=2294
      ("1000011100010011", "011"), -- i=2295
      ("1001011100010011", "011"), -- i=2296
      ("1010011100010011", "011"), -- i=2297
      ("1011011100010011", "011"), -- i=2298
      ("0100011100010000", "111"), -- i=2299
      ("1000011100010100", "100"), -- i=2300
      ("1001011100010100", "100"), -- i=2301
      ("1010011100010100", "100"), -- i=2302
      ("1011011100010100", "100"), -- i=2303
      ("0100011100010000", "111"), -- i=2304
      ("1000011100010101", "101"), -- i=2305
      ("1001011100010101", "101"), -- i=2306
      ("1010011100010101", "101"), -- i=2307
      ("1011011100010101", "101"), -- i=2308
      ("0100011100010000", "111"), -- i=2309
      ("1000011100010110", "110"), -- i=2310
      ("1001011100010110", "110"), -- i=2311
      ("1010011100010110", "110"), -- i=2312
      ("1011011100010110", "110"), -- i=2313
      ("0100011100010000", "111"), -- i=2314
      ("1000011100010111", "111"), -- i=2315
      ("1001011100010111", "111"), -- i=2316
      ("1010011100010111", "111"), -- i=2317
      ("1011011100010111", "111"), -- i=2318
      ("0100011100010000", "111"), -- i=2319
      ("1000011100100000", "000"), -- i=2320
      ("1001011100100000", "000"), -- i=2321
      ("1010011100100000", "000"), -- i=2322
      ("1011011100100000", "000"), -- i=2323
      ("0100011100100000", "111"), -- i=2324
      ("1000011100100001", "001"), -- i=2325
      ("1001011100100001", "001"), -- i=2326
      ("1010011100100001", "001"), -- i=2327
      ("1011011100100001", "001"), -- i=2328
      ("0100011100100000", "111"), -- i=2329
      ("1000011100100010", "010"), -- i=2330
      ("1001011100100010", "010"), -- i=2331
      ("1010011100100010", "010"), -- i=2332
      ("1011011100100010", "010"), -- i=2333
      ("0100011100100000", "111"), -- i=2334
      ("1000011100100011", "011"), -- i=2335
      ("1001011100100011", "011"), -- i=2336
      ("1010011100100011", "011"), -- i=2337
      ("1011011100100011", "011"), -- i=2338
      ("0100011100100000", "111"), -- i=2339
      ("1000011100100100", "100"), -- i=2340
      ("1001011100100100", "100"), -- i=2341
      ("1010011100100100", "100"), -- i=2342
      ("1011011100100100", "100"), -- i=2343
      ("0100011100100000", "111"), -- i=2344
      ("1000011100100101", "101"), -- i=2345
      ("1001011100100101", "101"), -- i=2346
      ("1010011100100101", "101"), -- i=2347
      ("1011011100100101", "101"), -- i=2348
      ("0100011100100000", "111"), -- i=2349
      ("1000011100100110", "110"), -- i=2350
      ("1001011100100110", "110"), -- i=2351
      ("1010011100100110", "110"), -- i=2352
      ("1011011100100110", "110"), -- i=2353
      ("0100011100100000", "111"), -- i=2354
      ("1000011100100111", "111"), -- i=2355
      ("1001011100100111", "111"), -- i=2356
      ("1010011100100111", "111"), -- i=2357
      ("1011011100100111", "111"), -- i=2358
      ("0100011100100000", "111"), -- i=2359
      ("1000011100110000", "000"), -- i=2360
      ("1001011100110000", "000"), -- i=2361
      ("1010011100110000", "000"), -- i=2362
      ("1011011100110000", "000"), -- i=2363
      ("0100011100110000", "111"), -- i=2364
      ("1000011100110001", "001"), -- i=2365
      ("1001011100110001", "001"), -- i=2366
      ("1010011100110001", "001"), -- i=2367
      ("1011011100110001", "001"), -- i=2368
      ("0100011100110000", "111"), -- i=2369
      ("1000011100110010", "010"), -- i=2370
      ("1001011100110010", "010"), -- i=2371
      ("1010011100110010", "010"), -- i=2372
      ("1011011100110010", "010"), -- i=2373
      ("0100011100110000", "111"), -- i=2374
      ("1000011100110011", "011"), -- i=2375
      ("1001011100110011", "011"), -- i=2376
      ("1010011100110011", "011"), -- i=2377
      ("1011011100110011", "011"), -- i=2378
      ("0100011100110000", "111"), -- i=2379
      ("1000011100110100", "100"), -- i=2380
      ("1001011100110100", "100"), -- i=2381
      ("1010011100110100", "100"), -- i=2382
      ("1011011100110100", "100"), -- i=2383
      ("0100011100110000", "111"), -- i=2384
      ("1000011100110101", "101"), -- i=2385
      ("1001011100110101", "101"), -- i=2386
      ("1010011100110101", "101"), -- i=2387
      ("1011011100110101", "101"), -- i=2388
      ("0100011100110000", "111"), -- i=2389
      ("1000011100110110", "110"), -- i=2390
      ("1001011100110110", "110"), -- i=2391
      ("1010011100110110", "110"), -- i=2392
      ("1011011100110110", "110"), -- i=2393
      ("0100011100110000", "111"), -- i=2394
      ("1000011100110111", "111"), -- i=2395
      ("1001011100110111", "111"), -- i=2396
      ("1010011100110111", "111"), -- i=2397
      ("1011011100110111", "111"), -- i=2398
      ("0100011100110000", "111"), -- i=2399
      ("1000011101000000", "000"), -- i=2400
      ("1001011101000000", "000"), -- i=2401
      ("1010011101000000", "000"), -- i=2402
      ("1011011101000000", "000"), -- i=2403
      ("0100011101000000", "111"), -- i=2404
      ("1000011101000001", "001"), -- i=2405
      ("1001011101000001", "001"), -- i=2406
      ("1010011101000001", "001"), -- i=2407
      ("1011011101000001", "001"), -- i=2408
      ("0100011101000000", "111"), -- i=2409
      ("1000011101000010", "010"), -- i=2410
      ("1001011101000010", "010"), -- i=2411
      ("1010011101000010", "010"), -- i=2412
      ("1011011101000010", "010"), -- i=2413
      ("0100011101000000", "111"), -- i=2414
      ("1000011101000011", "011"), -- i=2415
      ("1001011101000011", "011"), -- i=2416
      ("1010011101000011", "011"), -- i=2417
      ("1011011101000011", "011"), -- i=2418
      ("0100011101000000", "111"), -- i=2419
      ("1000011101000100", "100"), -- i=2420
      ("1001011101000100", "100"), -- i=2421
      ("1010011101000100", "100"), -- i=2422
      ("1011011101000100", "100"), -- i=2423
      ("0100011101000000", "111"), -- i=2424
      ("1000011101000101", "101"), -- i=2425
      ("1001011101000101", "101"), -- i=2426
      ("1010011101000101", "101"), -- i=2427
      ("1011011101000101", "101"), -- i=2428
      ("0100011101000000", "111"), -- i=2429
      ("1000011101000110", "110"), -- i=2430
      ("1001011101000110", "110"), -- i=2431
      ("1010011101000110", "110"), -- i=2432
      ("1011011101000110", "110"), -- i=2433
      ("0100011101000000", "111"), -- i=2434
      ("1000011101000111", "111"), -- i=2435
      ("1001011101000111", "111"), -- i=2436
      ("1010011101000111", "111"), -- i=2437
      ("1011011101000111", "111"), -- i=2438
      ("0100011101000000", "111"), -- i=2439
      ("1000011101010000", "000"), -- i=2440
      ("1001011101010000", "000"), -- i=2441
      ("1010011101010000", "000"), -- i=2442
      ("1011011101010000", "000"), -- i=2443
      ("0100011101010000", "111"), -- i=2444
      ("1000011101010001", "001"), -- i=2445
      ("1001011101010001", "001"), -- i=2446
      ("1010011101010001", "001"), -- i=2447
      ("1011011101010001", "001"), -- i=2448
      ("0100011101010000", "111"), -- i=2449
      ("1000011101010010", "010"), -- i=2450
      ("1001011101010010", "010"), -- i=2451
      ("1010011101010010", "010"), -- i=2452
      ("1011011101010010", "010"), -- i=2453
      ("0100011101010000", "111"), -- i=2454
      ("1000011101010011", "011"), -- i=2455
      ("1001011101010011", "011"), -- i=2456
      ("1010011101010011", "011"), -- i=2457
      ("1011011101010011", "011"), -- i=2458
      ("0100011101010000", "111"), -- i=2459
      ("1000011101010100", "100"), -- i=2460
      ("1001011101010100", "100"), -- i=2461
      ("1010011101010100", "100"), -- i=2462
      ("1011011101010100", "100"), -- i=2463
      ("0100011101010000", "111"), -- i=2464
      ("1000011101010101", "101"), -- i=2465
      ("1001011101010101", "101"), -- i=2466
      ("1010011101010101", "101"), -- i=2467
      ("1011011101010101", "101"), -- i=2468
      ("0100011101010000", "111"), -- i=2469
      ("1000011101010110", "110"), -- i=2470
      ("1001011101010110", "110"), -- i=2471
      ("1010011101010110", "110"), -- i=2472
      ("1011011101010110", "110"), -- i=2473
      ("0100011101010000", "111"), -- i=2474
      ("1000011101010111", "111"), -- i=2475
      ("1001011101010111", "111"), -- i=2476
      ("1010011101010111", "111"), -- i=2477
      ("1011011101010111", "111"), -- i=2478
      ("0100011101010000", "111"), -- i=2479
      ("1000011101100000", "000"), -- i=2480
      ("1001011101100000", "000"), -- i=2481
      ("1010011101100000", "000"), -- i=2482
      ("1011011101100000", "000"), -- i=2483
      ("0100011101100000", "111"), -- i=2484
      ("1000011101100001", "001"), -- i=2485
      ("1001011101100001", "001"), -- i=2486
      ("1010011101100001", "001"), -- i=2487
      ("1011011101100001", "001"), -- i=2488
      ("0100011101100000", "111"), -- i=2489
      ("1000011101100010", "010"), -- i=2490
      ("1001011101100010", "010"), -- i=2491
      ("1010011101100010", "010"), -- i=2492
      ("1011011101100010", "010"), -- i=2493
      ("0100011101100000", "111"), -- i=2494
      ("1000011101100011", "011"), -- i=2495
      ("1001011101100011", "011"), -- i=2496
      ("1010011101100011", "011"), -- i=2497
      ("1011011101100011", "011"), -- i=2498
      ("0100011101100000", "111"), -- i=2499
      ("1000011101100100", "100"), -- i=2500
      ("1001011101100100", "100"), -- i=2501
      ("1010011101100100", "100"), -- i=2502
      ("1011011101100100", "100"), -- i=2503
      ("0100011101100000", "111"), -- i=2504
      ("1000011101100101", "101"), -- i=2505
      ("1001011101100101", "101"), -- i=2506
      ("1010011101100101", "101"), -- i=2507
      ("1011011101100101", "101"), -- i=2508
      ("0100011101100000", "111"), -- i=2509
      ("1000011101100110", "110"), -- i=2510
      ("1001011101100110", "110"), -- i=2511
      ("1010011101100110", "110"), -- i=2512
      ("1011011101100110", "110"), -- i=2513
      ("0100011101100000", "111"), -- i=2514
      ("1000011101100111", "111"), -- i=2515
      ("1001011101100111", "111"), -- i=2516
      ("1010011101100111", "111"), -- i=2517
      ("1011011101100111", "111"), -- i=2518
      ("0100011101100000", "111"), -- i=2519
      ("1000011101110000", "000"), -- i=2520
      ("1001011101110000", "000"), -- i=2521
      ("1010011101110000", "000"), -- i=2522
      ("1011011101110000", "000"), -- i=2523
      ("0100011101110000", "111"), -- i=2524
      ("1000011101110001", "001"), -- i=2525
      ("1001011101110001", "001"), -- i=2526
      ("1010011101110001", "001"), -- i=2527
      ("1011011101110001", "001"), -- i=2528
      ("0100011101110000", "111"), -- i=2529
      ("1000011101110010", "010"), -- i=2530
      ("1001011101110010", "010"), -- i=2531
      ("1010011101110010", "010"), -- i=2532
      ("1011011101110010", "010"), -- i=2533
      ("0100011101110000", "111"), -- i=2534
      ("1000011101110011", "011"), -- i=2535
      ("1001011101110011", "011"), -- i=2536
      ("1010011101110011", "011"), -- i=2537
      ("1011011101110011", "011"), -- i=2538
      ("0100011101110000", "111"), -- i=2539
      ("1000011101110100", "100"), -- i=2540
      ("1001011101110100", "100"), -- i=2541
      ("1010011101110100", "100"), -- i=2542
      ("1011011101110100", "100"), -- i=2543
      ("0100011101110000", "111"), -- i=2544
      ("1000011101110101", "101"), -- i=2545
      ("1001011101110101", "101"), -- i=2546
      ("1010011101110101", "101"), -- i=2547
      ("1011011101110101", "101"), -- i=2548
      ("0100011101110000", "111"), -- i=2549
      ("1000011101110110", "110"), -- i=2550
      ("1001011101110110", "110"), -- i=2551
      ("1010011101110110", "110"), -- i=2552
      ("1011011101110110", "110"), -- i=2553
      ("0100011101110000", "111"), -- i=2554
      ("1000011101110111", "111"), -- i=2555
      ("1001011101110111", "111"), -- i=2556
      ("1010011101110111", "111"), -- i=2557
      ("1011011101110111", "111"), -- i=2558
      ("0100011101110000", "111"));
  begin
    for i in patterns'range loop
      INST <= patterns(i).INST;
      wait for 10 ns;
      assert std_match(ALUOP, patterns(i).ALUOP) OR (ALUOP = "ZZ" AND patterns(i).ALUOP = "ZZ")
        report "wrong value for ALUOP, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).ALUOP) & ", found " & to_string(ALUOP) severity error;assert std_match(RS1, patterns(i).RS1) OR (RS1 = "ZZZ" AND patterns(i).RS1 = "ZZZ")
        report "wrong value for RS1, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).RS1) & ", found " & to_string(RS1) severity error;assert std_match(RS2, patterns(i).RS2) OR (RS2 = "ZZZ" AND patterns(i).RS2 = "ZZZ")
        report "wrong value for RS2, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).RS2) & ", found " & to_string(RS2) severity error;assert std_match(WS, patterns(i).WS) OR (WS = "ZZZ" AND patterns(i).WS = "ZZZ")
        report "wrong value for WS, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).WS) & ", found " & to_string(WS) severity error;assert std_match(STR, patterns(i).STR) OR (STR = 'Z' AND patterns(i).STR = 'Z')
        report "wrong value for STR, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).STR) & ", found " & std_logic'image(STR) severity error;assert std_match(WE, patterns(i).WE) OR (WE = 'Z' AND patterns(i).WE = 'Z')
        report "wrong value for WE, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).WE) & ", found " & std_logic'image(WE) severity error;assert std_match(DMUX, patterns(i).DMUX) OR (DMUX = "ZZ" AND patterns(i).DMUX = "ZZ")
        report "wrong value for DMUX, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).DMUX) & ", found " & to_string(DMUX) severity error;assert std_match(LDR, patterns(i).LDR) OR (LDR = 'Z' AND patterns(i).LDR = 'Z')
        report "wrong value for LDR, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).LDR) & ", found " & std_logic'image(LDR) severity error;end loop;
    wait;
  end process;
end behav;
