//  A testbench for control_unit_STR_tb
`timescale 1us/1ns

module control_unit_STR_tb;
    reg [15:0] INST;
    wire [1:0] ALUOP;
    wire [2:0] RS1;
    wire [2:0] RS2;
    wire [2:0] WS;
    wire STR;
    wire WE;
    wire [1:0] DMUX;
    wire LDR;

  control_unit control_unit0 (
    .INST(INST),
    .ALUOP(ALUOP),
    .RS1(RS1),
    .RS2(RS2),
    .WS(WS),
    .STR(STR),
    .WE(WE),
    .DMUX(DMUX),
    .LDR(LDR)
  );

    reg [16:0] patterns[0:3583];
    integer i;

    initial begin
      patterns[0] = 17'b1000000000000000_0;
      patterns[1] = 17'b1001000000000000_0;
      patterns[2] = 17'b1010000000000000_0;
      patterns[3] = 17'b1011000000000000_0;
      patterns[4] = 17'b0101000000000000_0;
      patterns[5] = 17'b0100000000000000_1;
      patterns[6] = 17'b0000000001000010_0;
      patterns[7] = 17'b1000000000000001_0;
      patterns[8] = 17'b1001000000000001_0;
      patterns[9] = 17'b1010000000000001_0;
      patterns[10] = 17'b1011000000000001_0;
      patterns[11] = 17'b0101000000000000_0;
      patterns[12] = 17'b0100000000000000_1;
      patterns[13] = 17'b0000000011101000_0;
      patterns[14] = 17'b1000000000000010_0;
      patterns[15] = 17'b1001000000000010_0;
      patterns[16] = 17'b1010000000000010_0;
      patterns[17] = 17'b1011000000000010_0;
      patterns[18] = 17'b0101000000000000_0;
      patterns[19] = 17'b0100000000000000_1;
      patterns[20] = 17'b0000000001111000_0;
      patterns[21] = 17'b1000000000000011_0;
      patterns[22] = 17'b1001000000000011_0;
      patterns[23] = 17'b1010000000000011_0;
      patterns[24] = 17'b1011000000000011_0;
      patterns[25] = 17'b0101000000000000_0;
      patterns[26] = 17'b0100000000000000_1;
      patterns[27] = 17'b0000000001111001_0;
      patterns[28] = 17'b1000000000000100_0;
      patterns[29] = 17'b1001000000000100_0;
      patterns[30] = 17'b1010000000000100_0;
      patterns[31] = 17'b1011000000000100_0;
      patterns[32] = 17'b0101000000000000_0;
      patterns[33] = 17'b0100000000000000_1;
      patterns[34] = 17'b0000000000111011_0;
      patterns[35] = 17'b1000000000000101_0;
      patterns[36] = 17'b1001000000000101_0;
      patterns[37] = 17'b1010000000000101_0;
      patterns[38] = 17'b1011000000000101_0;
      patterns[39] = 17'b0101000000000000_0;
      patterns[40] = 17'b0100000000000000_1;
      patterns[41] = 17'b0000000010101110_0;
      patterns[42] = 17'b1000000000000110_0;
      patterns[43] = 17'b1001000000000110_0;
      patterns[44] = 17'b1010000000000110_0;
      patterns[45] = 17'b1011000000000110_0;
      patterns[46] = 17'b0101000000000000_0;
      patterns[47] = 17'b0100000000000000_1;
      patterns[48] = 17'b0000000010010010_0;
      patterns[49] = 17'b1000000000000111_0;
      patterns[50] = 17'b1001000000000111_0;
      patterns[51] = 17'b1010000000000111_0;
      patterns[52] = 17'b1011000000000111_0;
      patterns[53] = 17'b0101000000000000_0;
      patterns[54] = 17'b0100000000000000_1;
      patterns[55] = 17'b0000000010010110_0;
      patterns[56] = 17'b1000000000010000_0;
      patterns[57] = 17'b1001000000010000_0;
      patterns[58] = 17'b1010000000010000_0;
      patterns[59] = 17'b1011000000010000_0;
      patterns[60] = 17'b0101000000010000_0;
      patterns[61] = 17'b0100000000010000_1;
      patterns[62] = 17'b0000000000010001_0;
      patterns[63] = 17'b1000000000010001_0;
      patterns[64] = 17'b1001000000010001_0;
      patterns[65] = 17'b1010000000010001_0;
      patterns[66] = 17'b1011000000010001_0;
      patterns[67] = 17'b0101000000010000_0;
      patterns[68] = 17'b0100000000010000_1;
      patterns[69] = 17'b0000000010010001_0;
      patterns[70] = 17'b1000000000010010_0;
      patterns[71] = 17'b1001000000010010_0;
      patterns[72] = 17'b1010000000010010_0;
      patterns[73] = 17'b1011000000010010_0;
      patterns[74] = 17'b0101000000010000_0;
      patterns[75] = 17'b0100000000010000_1;
      patterns[76] = 17'b0000000011110100_0;
      patterns[77] = 17'b1000000000010011_0;
      patterns[78] = 17'b1001000000010011_0;
      patterns[79] = 17'b1010000000010011_0;
      patterns[80] = 17'b1011000000010011_0;
      patterns[81] = 17'b0101000000010000_0;
      patterns[82] = 17'b0100000000010000_1;
      patterns[83] = 17'b0000000000111111_0;
      patterns[84] = 17'b1000000000010100_0;
      patterns[85] = 17'b1001000000010100_0;
      patterns[86] = 17'b1010000000010100_0;
      patterns[87] = 17'b1011000000010100_0;
      patterns[88] = 17'b0101000000010000_0;
      patterns[89] = 17'b0100000000010000_1;
      patterns[90] = 17'b0000000000011100_0;
      patterns[91] = 17'b1000000000010101_0;
      patterns[92] = 17'b1001000000010101_0;
      patterns[93] = 17'b1010000000010101_0;
      patterns[94] = 17'b1011000000010101_0;
      patterns[95] = 17'b0101000000010000_0;
      patterns[96] = 17'b0100000000010000_1;
      patterns[97] = 17'b0000000001001111_0;
      patterns[98] = 17'b1000000000010110_0;
      patterns[99] = 17'b1001000000010110_0;
      patterns[100] = 17'b1010000000010110_0;
      patterns[101] = 17'b1011000000010110_0;
      patterns[102] = 17'b0101000000010000_0;
      patterns[103] = 17'b0100000000010000_1;
      patterns[104] = 17'b0000000010001010_0;
      patterns[105] = 17'b1000000000010111_0;
      patterns[106] = 17'b1001000000010111_0;
      patterns[107] = 17'b1010000000010111_0;
      patterns[108] = 17'b1011000000010111_0;
      patterns[109] = 17'b0101000000010000_0;
      patterns[110] = 17'b0100000000010000_1;
      patterns[111] = 17'b0000000001101111_0;
      patterns[112] = 17'b1000000000100000_0;
      patterns[113] = 17'b1001000000100000_0;
      patterns[114] = 17'b1010000000100000_0;
      patterns[115] = 17'b1011000000100000_0;
      patterns[116] = 17'b0101000000100000_0;
      patterns[117] = 17'b0100000000100000_1;
      patterns[118] = 17'b0000000010101101_0;
      patterns[119] = 17'b1000000000100001_0;
      patterns[120] = 17'b1001000000100001_0;
      patterns[121] = 17'b1010000000100001_0;
      patterns[122] = 17'b1011000000100001_0;
      patterns[123] = 17'b0101000000100000_0;
      patterns[124] = 17'b0100000000100000_1;
      patterns[125] = 17'b0000000010000100_0;
      patterns[126] = 17'b1000000000100010_0;
      patterns[127] = 17'b1001000000100010_0;
      patterns[128] = 17'b1010000000100010_0;
      patterns[129] = 17'b1011000000100010_0;
      patterns[130] = 17'b0101000000100000_0;
      patterns[131] = 17'b0100000000100000_1;
      patterns[132] = 17'b0000000011001001_0;
      patterns[133] = 17'b1000000000100011_0;
      patterns[134] = 17'b1001000000100011_0;
      patterns[135] = 17'b1010000000100011_0;
      patterns[136] = 17'b1011000000100011_0;
      patterns[137] = 17'b0101000000100000_0;
      patterns[138] = 17'b0100000000100000_1;
      patterns[139] = 17'b0000000010010111_0;
      patterns[140] = 17'b1000000000100100_0;
      patterns[141] = 17'b1001000000100100_0;
      patterns[142] = 17'b1010000000100100_0;
      patterns[143] = 17'b1011000000100100_0;
      patterns[144] = 17'b0101000000100000_0;
      patterns[145] = 17'b0100000000100000_1;
      patterns[146] = 17'b0000000001111001_0;
      patterns[147] = 17'b1000000000100101_0;
      patterns[148] = 17'b1001000000100101_0;
      patterns[149] = 17'b1010000000100101_0;
      patterns[150] = 17'b1011000000100101_0;
      patterns[151] = 17'b0101000000100000_0;
      patterns[152] = 17'b0100000000100000_1;
      patterns[153] = 17'b0000000000100101_0;
      patterns[154] = 17'b1000000000100110_0;
      patterns[155] = 17'b1001000000100110_0;
      patterns[156] = 17'b1010000000100110_0;
      patterns[157] = 17'b1011000000100110_0;
      patterns[158] = 17'b0101000000100000_0;
      patterns[159] = 17'b0100000000100000_1;
      patterns[160] = 17'b0000000000101110_0;
      patterns[161] = 17'b1000000000100111_0;
      patterns[162] = 17'b1001000000100111_0;
      patterns[163] = 17'b1010000000100111_0;
      patterns[164] = 17'b1011000000100111_0;
      patterns[165] = 17'b0101000000100000_0;
      patterns[166] = 17'b0100000000100000_1;
      patterns[167] = 17'b0000000010001001_0;
      patterns[168] = 17'b1000000000110000_0;
      patterns[169] = 17'b1001000000110000_0;
      patterns[170] = 17'b1010000000110000_0;
      patterns[171] = 17'b1011000000110000_0;
      patterns[172] = 17'b0101000000110000_0;
      patterns[173] = 17'b0100000000110000_1;
      patterns[174] = 17'b0000000011101110_0;
      patterns[175] = 17'b1000000000110001_0;
      patterns[176] = 17'b1001000000110001_0;
      patterns[177] = 17'b1010000000110001_0;
      patterns[178] = 17'b1011000000110001_0;
      patterns[179] = 17'b0101000000110000_0;
      patterns[180] = 17'b0100000000110000_1;
      patterns[181] = 17'b0000000001100011_0;
      patterns[182] = 17'b1000000000110010_0;
      patterns[183] = 17'b1001000000110010_0;
      patterns[184] = 17'b1010000000110010_0;
      patterns[185] = 17'b1011000000110010_0;
      patterns[186] = 17'b0101000000110000_0;
      patterns[187] = 17'b0100000000110000_1;
      patterns[188] = 17'b0000000011111101_0;
      patterns[189] = 17'b1000000000110011_0;
      patterns[190] = 17'b1001000000110011_0;
      patterns[191] = 17'b1010000000110011_0;
      patterns[192] = 17'b1011000000110011_0;
      patterns[193] = 17'b0101000000110000_0;
      patterns[194] = 17'b0100000000110000_1;
      patterns[195] = 17'b0000000010110100_0;
      patterns[196] = 17'b1000000000110100_0;
      patterns[197] = 17'b1001000000110100_0;
      patterns[198] = 17'b1010000000110100_0;
      patterns[199] = 17'b1011000000110100_0;
      patterns[200] = 17'b0101000000110000_0;
      patterns[201] = 17'b0100000000110000_1;
      patterns[202] = 17'b0000000011001010_0;
      patterns[203] = 17'b1000000000110101_0;
      patterns[204] = 17'b1001000000110101_0;
      patterns[205] = 17'b1010000000110101_0;
      patterns[206] = 17'b1011000000110101_0;
      patterns[207] = 17'b0101000000110000_0;
      patterns[208] = 17'b0100000000110000_1;
      patterns[209] = 17'b0000000000001001_0;
      patterns[210] = 17'b1000000000110110_0;
      patterns[211] = 17'b1001000000110110_0;
      patterns[212] = 17'b1010000000110110_0;
      patterns[213] = 17'b1011000000110110_0;
      patterns[214] = 17'b0101000000110000_0;
      patterns[215] = 17'b0100000000110000_1;
      patterns[216] = 17'b0000000000110001_0;
      patterns[217] = 17'b1000000000110111_0;
      patterns[218] = 17'b1001000000110111_0;
      patterns[219] = 17'b1010000000110111_0;
      patterns[220] = 17'b1011000000110111_0;
      patterns[221] = 17'b0101000000110000_0;
      patterns[222] = 17'b0100000000110000_1;
      patterns[223] = 17'b0000000011111011_0;
      patterns[224] = 17'b1000000001000000_0;
      patterns[225] = 17'b1001000001000000_0;
      patterns[226] = 17'b1010000001000000_0;
      patterns[227] = 17'b1011000001000000_0;
      patterns[228] = 17'b0101000001000000_0;
      patterns[229] = 17'b0100000001000000_1;
      patterns[230] = 17'b0000000011111011_0;
      patterns[231] = 17'b1000000001000001_0;
      patterns[232] = 17'b1001000001000001_0;
      patterns[233] = 17'b1010000001000001_0;
      patterns[234] = 17'b1011000001000001_0;
      patterns[235] = 17'b0101000001000000_0;
      patterns[236] = 17'b0100000001000000_1;
      patterns[237] = 17'b0000000011011110_0;
      patterns[238] = 17'b1000000001000010_0;
      patterns[239] = 17'b1001000001000010_0;
      patterns[240] = 17'b1010000001000010_0;
      patterns[241] = 17'b1011000001000010_0;
      patterns[242] = 17'b0101000001000000_0;
      patterns[243] = 17'b0100000001000000_1;
      patterns[244] = 17'b0000000001100001_0;
      patterns[245] = 17'b1000000001000011_0;
      patterns[246] = 17'b1001000001000011_0;
      patterns[247] = 17'b1010000001000011_0;
      patterns[248] = 17'b1011000001000011_0;
      patterns[249] = 17'b0101000001000000_0;
      patterns[250] = 17'b0100000001000000_1;
      patterns[251] = 17'b0000000011111100_0;
      patterns[252] = 17'b1000000001000100_0;
      patterns[253] = 17'b1001000001000100_0;
      patterns[254] = 17'b1010000001000100_0;
      patterns[255] = 17'b1011000001000100_0;
      patterns[256] = 17'b0101000001000000_0;
      patterns[257] = 17'b0100000001000000_1;
      patterns[258] = 17'b0000000000111001_0;
      patterns[259] = 17'b1000000001000101_0;
      patterns[260] = 17'b1001000001000101_0;
      patterns[261] = 17'b1010000001000101_0;
      patterns[262] = 17'b1011000001000101_0;
      patterns[263] = 17'b0101000001000000_0;
      patterns[264] = 17'b0100000001000000_1;
      patterns[265] = 17'b0000000000011100_0;
      patterns[266] = 17'b1000000001000110_0;
      patterns[267] = 17'b1001000001000110_0;
      patterns[268] = 17'b1010000001000110_0;
      patterns[269] = 17'b1011000001000110_0;
      patterns[270] = 17'b0101000001000000_0;
      patterns[271] = 17'b0100000001000000_1;
      patterns[272] = 17'b0000000010101000_0;
      patterns[273] = 17'b1000000001000111_0;
      patterns[274] = 17'b1001000001000111_0;
      patterns[275] = 17'b1010000001000111_0;
      patterns[276] = 17'b1011000001000111_0;
      patterns[277] = 17'b0101000001000000_0;
      patterns[278] = 17'b0100000001000000_1;
      patterns[279] = 17'b0000000001011100_0;
      patterns[280] = 17'b1000000001010000_0;
      patterns[281] = 17'b1001000001010000_0;
      patterns[282] = 17'b1010000001010000_0;
      patterns[283] = 17'b1011000001010000_0;
      patterns[284] = 17'b0101000001010000_0;
      patterns[285] = 17'b0100000001010000_1;
      patterns[286] = 17'b0000000011111110_0;
      patterns[287] = 17'b1000000001010001_0;
      patterns[288] = 17'b1001000001010001_0;
      patterns[289] = 17'b1010000001010001_0;
      patterns[290] = 17'b1011000001010001_0;
      patterns[291] = 17'b0101000001010000_0;
      patterns[292] = 17'b0100000001010000_1;
      patterns[293] = 17'b0000000010111001_0;
      patterns[294] = 17'b1000000001010010_0;
      patterns[295] = 17'b1001000001010010_0;
      patterns[296] = 17'b1010000001010010_0;
      patterns[297] = 17'b1011000001010010_0;
      patterns[298] = 17'b0101000001010000_0;
      patterns[299] = 17'b0100000001010000_1;
      patterns[300] = 17'b0000000000010100_0;
      patterns[301] = 17'b1000000001010011_0;
      patterns[302] = 17'b1001000001010011_0;
      patterns[303] = 17'b1010000001010011_0;
      patterns[304] = 17'b1011000001010011_0;
      patterns[305] = 17'b0101000001010000_0;
      patterns[306] = 17'b0100000001010000_1;
      patterns[307] = 17'b0000000001011000_0;
      patterns[308] = 17'b1000000001010100_0;
      patterns[309] = 17'b1001000001010100_0;
      patterns[310] = 17'b1010000001010100_0;
      patterns[311] = 17'b1011000001010100_0;
      patterns[312] = 17'b0101000001010000_0;
      patterns[313] = 17'b0100000001010000_1;
      patterns[314] = 17'b0000000010010100_0;
      patterns[315] = 17'b1000000001010101_0;
      patterns[316] = 17'b1001000001010101_0;
      patterns[317] = 17'b1010000001010101_0;
      patterns[318] = 17'b1011000001010101_0;
      patterns[319] = 17'b0101000001010000_0;
      patterns[320] = 17'b0100000001010000_1;
      patterns[321] = 17'b0000000010101111_0;
      patterns[322] = 17'b1000000001010110_0;
      patterns[323] = 17'b1001000001010110_0;
      patterns[324] = 17'b1010000001010110_0;
      patterns[325] = 17'b1011000001010110_0;
      patterns[326] = 17'b0101000001010000_0;
      patterns[327] = 17'b0100000001010000_1;
      patterns[328] = 17'b0000000011010100_0;
      patterns[329] = 17'b1000000001010111_0;
      patterns[330] = 17'b1001000001010111_0;
      patterns[331] = 17'b1010000001010111_0;
      patterns[332] = 17'b1011000001010111_0;
      patterns[333] = 17'b0101000001010000_0;
      patterns[334] = 17'b0100000001010000_1;
      patterns[335] = 17'b0000000010110001_0;
      patterns[336] = 17'b1000000001100000_0;
      patterns[337] = 17'b1001000001100000_0;
      patterns[338] = 17'b1010000001100000_0;
      patterns[339] = 17'b1011000001100000_0;
      patterns[340] = 17'b0101000001100000_0;
      patterns[341] = 17'b0100000001100000_1;
      patterns[342] = 17'b0000000010011110_0;
      patterns[343] = 17'b1000000001100001_0;
      patterns[344] = 17'b1001000001100001_0;
      patterns[345] = 17'b1010000001100001_0;
      patterns[346] = 17'b1011000001100001_0;
      patterns[347] = 17'b0101000001100000_0;
      patterns[348] = 17'b0100000001100000_1;
      patterns[349] = 17'b0000000000110110_0;
      patterns[350] = 17'b1000000001100010_0;
      patterns[351] = 17'b1001000001100010_0;
      patterns[352] = 17'b1010000001100010_0;
      patterns[353] = 17'b1011000001100010_0;
      patterns[354] = 17'b0101000001100000_0;
      patterns[355] = 17'b0100000001100000_1;
      patterns[356] = 17'b0000000010000111_0;
      patterns[357] = 17'b1000000001100011_0;
      patterns[358] = 17'b1001000001100011_0;
      patterns[359] = 17'b1010000001100011_0;
      patterns[360] = 17'b1011000001100011_0;
      patterns[361] = 17'b0101000001100000_0;
      patterns[362] = 17'b0100000001100000_1;
      patterns[363] = 17'b0000000010100000_0;
      patterns[364] = 17'b1000000001100100_0;
      patterns[365] = 17'b1001000001100100_0;
      patterns[366] = 17'b1010000001100100_0;
      patterns[367] = 17'b1011000001100100_0;
      patterns[368] = 17'b0101000001100000_0;
      patterns[369] = 17'b0100000001100000_1;
      patterns[370] = 17'b0000000000101000_0;
      patterns[371] = 17'b1000000001100101_0;
      patterns[372] = 17'b1001000001100101_0;
      patterns[373] = 17'b1010000001100101_0;
      patterns[374] = 17'b1011000001100101_0;
      patterns[375] = 17'b0101000001100000_0;
      patterns[376] = 17'b0100000001100000_1;
      patterns[377] = 17'b0000000010000111_0;
      patterns[378] = 17'b1000000001100110_0;
      patterns[379] = 17'b1001000001100110_0;
      patterns[380] = 17'b1010000001100110_0;
      patterns[381] = 17'b1011000001100110_0;
      patterns[382] = 17'b0101000001100000_0;
      patterns[383] = 17'b0100000001100000_1;
      patterns[384] = 17'b0000000001001110_0;
      patterns[385] = 17'b1000000001100111_0;
      patterns[386] = 17'b1001000001100111_0;
      patterns[387] = 17'b1010000001100111_0;
      patterns[388] = 17'b1011000001100111_0;
      patterns[389] = 17'b0101000001100000_0;
      patterns[390] = 17'b0100000001100000_1;
      patterns[391] = 17'b0000000010001101_0;
      patterns[392] = 17'b1000000001110000_0;
      patterns[393] = 17'b1001000001110000_0;
      patterns[394] = 17'b1010000001110000_0;
      patterns[395] = 17'b1011000001110000_0;
      patterns[396] = 17'b0101000001110000_0;
      patterns[397] = 17'b0100000001110000_1;
      patterns[398] = 17'b0000000010011010_0;
      patterns[399] = 17'b1000000001110001_0;
      patterns[400] = 17'b1001000001110001_0;
      patterns[401] = 17'b1010000001110001_0;
      patterns[402] = 17'b1011000001110001_0;
      patterns[403] = 17'b0101000001110000_0;
      patterns[404] = 17'b0100000001110000_1;
      patterns[405] = 17'b0000000001011001_0;
      patterns[406] = 17'b1000000001110010_0;
      patterns[407] = 17'b1001000001110010_0;
      patterns[408] = 17'b1010000001110010_0;
      patterns[409] = 17'b1011000001110010_0;
      patterns[410] = 17'b0101000001110000_0;
      patterns[411] = 17'b0100000001110000_1;
      patterns[412] = 17'b0000000011010111_0;
      patterns[413] = 17'b1000000001110011_0;
      patterns[414] = 17'b1001000001110011_0;
      patterns[415] = 17'b1010000001110011_0;
      patterns[416] = 17'b1011000001110011_0;
      patterns[417] = 17'b0101000001110000_0;
      patterns[418] = 17'b0100000001110000_1;
      patterns[419] = 17'b0000000011010011_0;
      patterns[420] = 17'b1000000001110100_0;
      patterns[421] = 17'b1001000001110100_0;
      patterns[422] = 17'b1010000001110100_0;
      patterns[423] = 17'b1011000001110100_0;
      patterns[424] = 17'b0101000001110000_0;
      patterns[425] = 17'b0100000001110000_1;
      patterns[426] = 17'b0000000000000000_0;
      patterns[427] = 17'b1000000001110101_0;
      patterns[428] = 17'b1001000001110101_0;
      patterns[429] = 17'b1010000001110101_0;
      patterns[430] = 17'b1011000001110101_0;
      patterns[431] = 17'b0101000001110000_0;
      patterns[432] = 17'b0100000001110000_1;
      patterns[433] = 17'b0000000000100011_0;
      patterns[434] = 17'b1000000001110110_0;
      patterns[435] = 17'b1001000001110110_0;
      patterns[436] = 17'b1010000001110110_0;
      patterns[437] = 17'b1011000001110110_0;
      patterns[438] = 17'b0101000001110000_0;
      patterns[439] = 17'b0100000001110000_1;
      patterns[440] = 17'b0000000010100001_0;
      patterns[441] = 17'b1000000001110111_0;
      patterns[442] = 17'b1001000001110111_0;
      patterns[443] = 17'b1010000001110111_0;
      patterns[444] = 17'b1011000001110111_0;
      patterns[445] = 17'b0101000001110000_0;
      patterns[446] = 17'b0100000001110000_1;
      patterns[447] = 17'b0000000000001010_0;
      patterns[448] = 17'b1000000100000000_0;
      patterns[449] = 17'b1001000100000000_0;
      patterns[450] = 17'b1010000100000000_0;
      patterns[451] = 17'b1011000100000000_0;
      patterns[452] = 17'b0101000100000000_0;
      patterns[453] = 17'b0100000100000000_1;
      patterns[454] = 17'b0000000100011100_0;
      patterns[455] = 17'b1000000100000001_0;
      patterns[456] = 17'b1001000100000001_0;
      patterns[457] = 17'b1010000100000001_0;
      patterns[458] = 17'b1011000100000001_0;
      patterns[459] = 17'b0101000100000000_0;
      patterns[460] = 17'b0100000100000000_1;
      patterns[461] = 17'b0000000111100001_0;
      patterns[462] = 17'b1000000100000010_0;
      patterns[463] = 17'b1001000100000010_0;
      patterns[464] = 17'b1010000100000010_0;
      patterns[465] = 17'b1011000100000010_0;
      patterns[466] = 17'b0101000100000000_0;
      patterns[467] = 17'b0100000100000000_1;
      patterns[468] = 17'b0000000110110011_0;
      patterns[469] = 17'b1000000100000011_0;
      patterns[470] = 17'b1001000100000011_0;
      patterns[471] = 17'b1010000100000011_0;
      patterns[472] = 17'b1011000100000011_0;
      patterns[473] = 17'b0101000100000000_0;
      patterns[474] = 17'b0100000100000000_1;
      patterns[475] = 17'b0000000111010111_0;
      patterns[476] = 17'b1000000100000100_0;
      patterns[477] = 17'b1001000100000100_0;
      patterns[478] = 17'b1010000100000100_0;
      patterns[479] = 17'b1011000100000100_0;
      patterns[480] = 17'b0101000100000000_0;
      patterns[481] = 17'b0100000100000000_1;
      patterns[482] = 17'b0000000101000011_0;
      patterns[483] = 17'b1000000100000101_0;
      patterns[484] = 17'b1001000100000101_0;
      patterns[485] = 17'b1010000100000101_0;
      patterns[486] = 17'b1011000100000101_0;
      patterns[487] = 17'b0101000100000000_0;
      patterns[488] = 17'b0100000100000000_1;
      patterns[489] = 17'b0000000111011010_0;
      patterns[490] = 17'b1000000100000110_0;
      patterns[491] = 17'b1001000100000110_0;
      patterns[492] = 17'b1010000100000110_0;
      patterns[493] = 17'b1011000100000110_0;
      patterns[494] = 17'b0101000100000000_0;
      patterns[495] = 17'b0100000100000000_1;
      patterns[496] = 17'b0000000110011100_0;
      patterns[497] = 17'b1000000100000111_0;
      patterns[498] = 17'b1001000100000111_0;
      patterns[499] = 17'b1010000100000111_0;
      patterns[500] = 17'b1011000100000111_0;
      patterns[501] = 17'b0101000100000000_0;
      patterns[502] = 17'b0100000100000000_1;
      patterns[503] = 17'b0000000110011000_0;
      patterns[504] = 17'b1000000100010000_0;
      patterns[505] = 17'b1001000100010000_0;
      patterns[506] = 17'b1010000100010000_0;
      patterns[507] = 17'b1011000100010000_0;
      patterns[508] = 17'b0101000100010000_0;
      patterns[509] = 17'b0100000100010000_1;
      patterns[510] = 17'b0000000110100001_0;
      patterns[511] = 17'b1000000100010001_0;
      patterns[512] = 17'b1001000100010001_0;
      patterns[513] = 17'b1010000100010001_0;
      patterns[514] = 17'b1011000100010001_0;
      patterns[515] = 17'b0101000100010000_0;
      patterns[516] = 17'b0100000100010000_1;
      patterns[517] = 17'b0000000111011010_0;
      patterns[518] = 17'b1000000100010010_0;
      patterns[519] = 17'b1001000100010010_0;
      patterns[520] = 17'b1010000100010010_0;
      patterns[521] = 17'b1011000100010010_0;
      patterns[522] = 17'b0101000100010000_0;
      patterns[523] = 17'b0100000100010000_1;
      patterns[524] = 17'b0000000100111100_0;
      patterns[525] = 17'b1000000100010011_0;
      patterns[526] = 17'b1001000100010011_0;
      patterns[527] = 17'b1010000100010011_0;
      patterns[528] = 17'b1011000100010011_0;
      patterns[529] = 17'b0101000100010000_0;
      patterns[530] = 17'b0100000100010000_1;
      patterns[531] = 17'b0000000111011000_0;
      patterns[532] = 17'b1000000100010100_0;
      patterns[533] = 17'b1001000100010100_0;
      patterns[534] = 17'b1010000100010100_0;
      patterns[535] = 17'b1011000100010100_0;
      patterns[536] = 17'b0101000100010000_0;
      patterns[537] = 17'b0100000100010000_1;
      patterns[538] = 17'b0000000110101011_0;
      patterns[539] = 17'b1000000100010101_0;
      patterns[540] = 17'b1001000100010101_0;
      patterns[541] = 17'b1010000100010101_0;
      patterns[542] = 17'b1011000100010101_0;
      patterns[543] = 17'b0101000100010000_0;
      patterns[544] = 17'b0100000100010000_1;
      patterns[545] = 17'b0000000111111000_0;
      patterns[546] = 17'b1000000100010110_0;
      patterns[547] = 17'b1001000100010110_0;
      patterns[548] = 17'b1010000100010110_0;
      patterns[549] = 17'b1011000100010110_0;
      patterns[550] = 17'b0101000100010000_0;
      patterns[551] = 17'b0100000100010000_1;
      patterns[552] = 17'b0000000111011110_0;
      patterns[553] = 17'b1000000100010111_0;
      patterns[554] = 17'b1001000100010111_0;
      patterns[555] = 17'b1010000100010111_0;
      patterns[556] = 17'b1011000100010111_0;
      patterns[557] = 17'b0101000100010000_0;
      patterns[558] = 17'b0100000100010000_1;
      patterns[559] = 17'b0000000111000100_0;
      patterns[560] = 17'b1000000100100000_0;
      patterns[561] = 17'b1001000100100000_0;
      patterns[562] = 17'b1010000100100000_0;
      patterns[563] = 17'b1011000100100000_0;
      patterns[564] = 17'b0101000100100000_0;
      patterns[565] = 17'b0100000100100000_1;
      patterns[566] = 17'b0000000110001101_0;
      patterns[567] = 17'b1000000100100001_0;
      patterns[568] = 17'b1001000100100001_0;
      patterns[569] = 17'b1010000100100001_0;
      patterns[570] = 17'b1011000100100001_0;
      patterns[571] = 17'b0101000100100000_0;
      patterns[572] = 17'b0100000100100000_1;
      patterns[573] = 17'b0000000100011101_0;
      patterns[574] = 17'b1000000100100010_0;
      patterns[575] = 17'b1001000100100010_0;
      patterns[576] = 17'b1010000100100010_0;
      patterns[577] = 17'b1011000100100010_0;
      patterns[578] = 17'b0101000100100000_0;
      patterns[579] = 17'b0100000100100000_1;
      patterns[580] = 17'b0000000101110110_0;
      patterns[581] = 17'b1000000100100011_0;
      patterns[582] = 17'b1001000100100011_0;
      patterns[583] = 17'b1010000100100011_0;
      patterns[584] = 17'b1011000100100011_0;
      patterns[585] = 17'b0101000100100000_0;
      patterns[586] = 17'b0100000100100000_1;
      patterns[587] = 17'b0000000110011110_0;
      patterns[588] = 17'b1000000100100100_0;
      patterns[589] = 17'b1001000100100100_0;
      patterns[590] = 17'b1010000100100100_0;
      patterns[591] = 17'b1011000100100100_0;
      patterns[592] = 17'b0101000100100000_0;
      patterns[593] = 17'b0100000100100000_1;
      patterns[594] = 17'b0000000101001001_0;
      patterns[595] = 17'b1000000100100101_0;
      patterns[596] = 17'b1001000100100101_0;
      patterns[597] = 17'b1010000100100101_0;
      patterns[598] = 17'b1011000100100101_0;
      patterns[599] = 17'b0101000100100000_0;
      patterns[600] = 17'b0100000100100000_1;
      patterns[601] = 17'b0000000100111011_0;
      patterns[602] = 17'b1000000100100110_0;
      patterns[603] = 17'b1001000100100110_0;
      patterns[604] = 17'b1010000100100110_0;
      patterns[605] = 17'b1011000100100110_0;
      patterns[606] = 17'b0101000100100000_0;
      patterns[607] = 17'b0100000100100000_1;
      patterns[608] = 17'b0000000101101111_0;
      patterns[609] = 17'b1000000100100111_0;
      patterns[610] = 17'b1001000100100111_0;
      patterns[611] = 17'b1010000100100111_0;
      patterns[612] = 17'b1011000100100111_0;
      patterns[613] = 17'b0101000100100000_0;
      patterns[614] = 17'b0100000100100000_1;
      patterns[615] = 17'b0000000101111010_0;
      patterns[616] = 17'b1000000100110000_0;
      patterns[617] = 17'b1001000100110000_0;
      patterns[618] = 17'b1010000100110000_0;
      patterns[619] = 17'b1011000100110000_0;
      patterns[620] = 17'b0101000100110000_0;
      patterns[621] = 17'b0100000100110000_1;
      patterns[622] = 17'b0000000110111010_0;
      patterns[623] = 17'b1000000100110001_0;
      patterns[624] = 17'b1001000100110001_0;
      patterns[625] = 17'b1010000100110001_0;
      patterns[626] = 17'b1011000100110001_0;
      patterns[627] = 17'b0101000100110000_0;
      patterns[628] = 17'b0100000100110000_1;
      patterns[629] = 17'b0000000100110010_0;
      patterns[630] = 17'b1000000100110010_0;
      patterns[631] = 17'b1001000100110010_0;
      patterns[632] = 17'b1010000100110010_0;
      patterns[633] = 17'b1011000100110010_0;
      patterns[634] = 17'b0101000100110000_0;
      patterns[635] = 17'b0100000100110000_1;
      patterns[636] = 17'b0000000101000110_0;
      patterns[637] = 17'b1000000100110011_0;
      patterns[638] = 17'b1001000100110011_0;
      patterns[639] = 17'b1010000100110011_0;
      patterns[640] = 17'b1011000100110011_0;
      patterns[641] = 17'b0101000100110000_0;
      patterns[642] = 17'b0100000100110000_1;
      patterns[643] = 17'b0000000101100010_0;
      patterns[644] = 17'b1000000100110100_0;
      patterns[645] = 17'b1001000100110100_0;
      patterns[646] = 17'b1010000100110100_0;
      patterns[647] = 17'b1011000100110100_0;
      patterns[648] = 17'b0101000100110000_0;
      patterns[649] = 17'b0100000100110000_1;
      patterns[650] = 17'b0000000100010010_0;
      patterns[651] = 17'b1000000100110101_0;
      patterns[652] = 17'b1001000100110101_0;
      patterns[653] = 17'b1010000100110101_0;
      patterns[654] = 17'b1011000100110101_0;
      patterns[655] = 17'b0101000100110000_0;
      patterns[656] = 17'b0100000100110000_1;
      patterns[657] = 17'b0000000101010001_0;
      patterns[658] = 17'b1000000100110110_0;
      patterns[659] = 17'b1001000100110110_0;
      patterns[660] = 17'b1010000100110110_0;
      patterns[661] = 17'b1011000100110110_0;
      patterns[662] = 17'b0101000100110000_0;
      patterns[663] = 17'b0100000100110000_1;
      patterns[664] = 17'b0000000101101000_0;
      patterns[665] = 17'b1000000100110111_0;
      patterns[666] = 17'b1001000100110111_0;
      patterns[667] = 17'b1010000100110111_0;
      patterns[668] = 17'b1011000100110111_0;
      patterns[669] = 17'b0101000100110000_0;
      patterns[670] = 17'b0100000100110000_1;
      patterns[671] = 17'b0000000101100101_0;
      patterns[672] = 17'b1000000101000000_0;
      patterns[673] = 17'b1001000101000000_0;
      patterns[674] = 17'b1010000101000000_0;
      patterns[675] = 17'b1011000101000000_0;
      patterns[676] = 17'b0101000101000000_0;
      patterns[677] = 17'b0100000101000000_1;
      patterns[678] = 17'b0000000110110001_0;
      patterns[679] = 17'b1000000101000001_0;
      patterns[680] = 17'b1001000101000001_0;
      patterns[681] = 17'b1010000101000001_0;
      patterns[682] = 17'b1011000101000001_0;
      patterns[683] = 17'b0101000101000000_0;
      patterns[684] = 17'b0100000101000000_1;
      patterns[685] = 17'b0000000101100001_0;
      patterns[686] = 17'b1000000101000010_0;
      patterns[687] = 17'b1001000101000010_0;
      patterns[688] = 17'b1010000101000010_0;
      patterns[689] = 17'b1011000101000010_0;
      patterns[690] = 17'b0101000101000000_0;
      patterns[691] = 17'b0100000101000000_1;
      patterns[692] = 17'b0000000100010111_0;
      patterns[693] = 17'b1000000101000011_0;
      patterns[694] = 17'b1001000101000011_0;
      patterns[695] = 17'b1010000101000011_0;
      patterns[696] = 17'b1011000101000011_0;
      patterns[697] = 17'b0101000101000000_0;
      patterns[698] = 17'b0100000101000000_1;
      patterns[699] = 17'b0000000111110100_0;
      patterns[700] = 17'b1000000101000100_0;
      patterns[701] = 17'b1001000101000100_0;
      patterns[702] = 17'b1010000101000100_0;
      patterns[703] = 17'b1011000101000100_0;
      patterns[704] = 17'b0101000101000000_0;
      patterns[705] = 17'b0100000101000000_1;
      patterns[706] = 17'b0000000111101101_0;
      patterns[707] = 17'b1000000101000101_0;
      patterns[708] = 17'b1001000101000101_0;
      patterns[709] = 17'b1010000101000101_0;
      patterns[710] = 17'b1011000101000101_0;
      patterns[711] = 17'b0101000101000000_0;
      patterns[712] = 17'b0100000101000000_1;
      patterns[713] = 17'b0000000100111001_0;
      patterns[714] = 17'b1000000101000110_0;
      patterns[715] = 17'b1001000101000110_0;
      patterns[716] = 17'b1010000101000110_0;
      patterns[717] = 17'b1011000101000110_0;
      patterns[718] = 17'b0101000101000000_0;
      patterns[719] = 17'b0100000101000000_1;
      patterns[720] = 17'b0000000111110100_0;
      patterns[721] = 17'b1000000101000111_0;
      patterns[722] = 17'b1001000101000111_0;
      patterns[723] = 17'b1010000101000111_0;
      patterns[724] = 17'b1011000101000111_0;
      patterns[725] = 17'b0101000101000000_0;
      patterns[726] = 17'b0100000101000000_1;
      patterns[727] = 17'b0000000101100001_0;
      patterns[728] = 17'b1000000101010000_0;
      patterns[729] = 17'b1001000101010000_0;
      patterns[730] = 17'b1010000101010000_0;
      patterns[731] = 17'b1011000101010000_0;
      patterns[732] = 17'b0101000101010000_0;
      patterns[733] = 17'b0100000101010000_1;
      patterns[734] = 17'b0000000101010011_0;
      patterns[735] = 17'b1000000101010001_0;
      patterns[736] = 17'b1001000101010001_0;
      patterns[737] = 17'b1010000101010001_0;
      patterns[738] = 17'b1011000101010001_0;
      patterns[739] = 17'b0101000101010000_0;
      patterns[740] = 17'b0100000101010000_1;
      patterns[741] = 17'b0000000111101000_0;
      patterns[742] = 17'b1000000101010010_0;
      patterns[743] = 17'b1001000101010010_0;
      patterns[744] = 17'b1010000101010010_0;
      patterns[745] = 17'b1011000101010010_0;
      patterns[746] = 17'b0101000101010000_0;
      patterns[747] = 17'b0100000101010000_1;
      patterns[748] = 17'b0000000110011011_0;
      patterns[749] = 17'b1000000101010011_0;
      patterns[750] = 17'b1001000101010011_0;
      patterns[751] = 17'b1010000101010011_0;
      patterns[752] = 17'b1011000101010011_0;
      patterns[753] = 17'b0101000101010000_0;
      patterns[754] = 17'b0100000101010000_1;
      patterns[755] = 17'b0000000101001000_0;
      patterns[756] = 17'b1000000101010100_0;
      patterns[757] = 17'b1001000101010100_0;
      patterns[758] = 17'b1010000101010100_0;
      patterns[759] = 17'b1011000101010100_0;
      patterns[760] = 17'b0101000101010000_0;
      patterns[761] = 17'b0100000101010000_1;
      patterns[762] = 17'b0000000101000000_0;
      patterns[763] = 17'b1000000101010101_0;
      patterns[764] = 17'b1001000101010101_0;
      patterns[765] = 17'b1010000101010101_0;
      patterns[766] = 17'b1011000101010101_0;
      patterns[767] = 17'b0101000101010000_0;
      patterns[768] = 17'b0100000101010000_1;
      patterns[769] = 17'b0000000110100000_0;
      patterns[770] = 17'b1000000101010110_0;
      patterns[771] = 17'b1001000101010110_0;
      patterns[772] = 17'b1010000101010110_0;
      patterns[773] = 17'b1011000101010110_0;
      patterns[774] = 17'b0101000101010000_0;
      patterns[775] = 17'b0100000101010000_1;
      patterns[776] = 17'b0000000100110101_0;
      patterns[777] = 17'b1000000101010111_0;
      patterns[778] = 17'b1001000101010111_0;
      patterns[779] = 17'b1010000101010111_0;
      patterns[780] = 17'b1011000101010111_0;
      patterns[781] = 17'b0101000101010000_0;
      patterns[782] = 17'b0100000101010000_1;
      patterns[783] = 17'b0000000100110011_0;
      patterns[784] = 17'b1000000101100000_0;
      patterns[785] = 17'b1001000101100000_0;
      patterns[786] = 17'b1010000101100000_0;
      patterns[787] = 17'b1011000101100000_0;
      patterns[788] = 17'b0101000101100000_0;
      patterns[789] = 17'b0100000101100000_1;
      patterns[790] = 17'b0000000100001111_0;
      patterns[791] = 17'b1000000101100001_0;
      patterns[792] = 17'b1001000101100001_0;
      patterns[793] = 17'b1010000101100001_0;
      patterns[794] = 17'b1011000101100001_0;
      patterns[795] = 17'b0101000101100000_0;
      patterns[796] = 17'b0100000101100000_1;
      patterns[797] = 17'b0000000110100001_0;
      patterns[798] = 17'b1000000101100010_0;
      patterns[799] = 17'b1001000101100010_0;
      patterns[800] = 17'b1010000101100010_0;
      patterns[801] = 17'b1011000101100010_0;
      patterns[802] = 17'b0101000101100000_0;
      patterns[803] = 17'b0100000101100000_1;
      patterns[804] = 17'b0000000101000101_0;
      patterns[805] = 17'b1000000101100011_0;
      patterns[806] = 17'b1001000101100011_0;
      patterns[807] = 17'b1010000101100011_0;
      patterns[808] = 17'b1011000101100011_0;
      patterns[809] = 17'b0101000101100000_0;
      patterns[810] = 17'b0100000101100000_1;
      patterns[811] = 17'b0000000110110111_0;
      patterns[812] = 17'b1000000101100100_0;
      patterns[813] = 17'b1001000101100100_0;
      patterns[814] = 17'b1010000101100100_0;
      patterns[815] = 17'b1011000101100100_0;
      patterns[816] = 17'b0101000101100000_0;
      patterns[817] = 17'b0100000101100000_1;
      patterns[818] = 17'b0000000100101001_0;
      patterns[819] = 17'b1000000101100101_0;
      patterns[820] = 17'b1001000101100101_0;
      patterns[821] = 17'b1010000101100101_0;
      patterns[822] = 17'b1011000101100101_0;
      patterns[823] = 17'b0101000101100000_0;
      patterns[824] = 17'b0100000101100000_1;
      patterns[825] = 17'b0000000110101100_0;
      patterns[826] = 17'b1000000101100110_0;
      patterns[827] = 17'b1001000101100110_0;
      patterns[828] = 17'b1010000101100110_0;
      patterns[829] = 17'b1011000101100110_0;
      patterns[830] = 17'b0101000101100000_0;
      patterns[831] = 17'b0100000101100000_1;
      patterns[832] = 17'b0000000111011000_0;
      patterns[833] = 17'b1000000101100111_0;
      patterns[834] = 17'b1001000101100111_0;
      patterns[835] = 17'b1010000101100111_0;
      patterns[836] = 17'b1011000101100111_0;
      patterns[837] = 17'b0101000101100000_0;
      patterns[838] = 17'b0100000101100000_1;
      patterns[839] = 17'b0000000111111011_0;
      patterns[840] = 17'b1000000101110000_0;
      patterns[841] = 17'b1001000101110000_0;
      patterns[842] = 17'b1010000101110000_0;
      patterns[843] = 17'b1011000101110000_0;
      patterns[844] = 17'b0101000101110000_0;
      patterns[845] = 17'b0100000101110000_1;
      patterns[846] = 17'b0000000100000110_0;
      patterns[847] = 17'b1000000101110001_0;
      patterns[848] = 17'b1001000101110001_0;
      patterns[849] = 17'b1010000101110001_0;
      patterns[850] = 17'b1011000101110001_0;
      patterns[851] = 17'b0101000101110000_0;
      patterns[852] = 17'b0100000101110000_1;
      patterns[853] = 17'b0000000110001110_0;
      patterns[854] = 17'b1000000101110010_0;
      patterns[855] = 17'b1001000101110010_0;
      patterns[856] = 17'b1010000101110010_0;
      patterns[857] = 17'b1011000101110010_0;
      patterns[858] = 17'b0101000101110000_0;
      patterns[859] = 17'b0100000101110000_1;
      patterns[860] = 17'b0000000101110100_0;
      patterns[861] = 17'b1000000101110011_0;
      patterns[862] = 17'b1001000101110011_0;
      patterns[863] = 17'b1010000101110011_0;
      patterns[864] = 17'b1011000101110011_0;
      patterns[865] = 17'b0101000101110000_0;
      patterns[866] = 17'b0100000101110000_1;
      patterns[867] = 17'b0000000110001000_0;
      patterns[868] = 17'b1000000101110100_0;
      patterns[869] = 17'b1001000101110100_0;
      patterns[870] = 17'b1010000101110100_0;
      patterns[871] = 17'b1011000101110100_0;
      patterns[872] = 17'b0101000101110000_0;
      patterns[873] = 17'b0100000101110000_1;
      patterns[874] = 17'b0000000111101111_0;
      patterns[875] = 17'b1000000101110101_0;
      patterns[876] = 17'b1001000101110101_0;
      patterns[877] = 17'b1010000101110101_0;
      patterns[878] = 17'b1011000101110101_0;
      patterns[879] = 17'b0101000101110000_0;
      patterns[880] = 17'b0100000101110000_1;
      patterns[881] = 17'b0000000110111110_0;
      patterns[882] = 17'b1000000101110110_0;
      patterns[883] = 17'b1001000101110110_0;
      patterns[884] = 17'b1010000101110110_0;
      patterns[885] = 17'b1011000101110110_0;
      patterns[886] = 17'b0101000101110000_0;
      patterns[887] = 17'b0100000101110000_1;
      patterns[888] = 17'b0000000101010111_0;
      patterns[889] = 17'b1000000101110111_0;
      patterns[890] = 17'b1001000101110111_0;
      patterns[891] = 17'b1010000101110111_0;
      patterns[892] = 17'b1011000101110111_0;
      patterns[893] = 17'b0101000101110000_0;
      patterns[894] = 17'b0100000101110000_1;
      patterns[895] = 17'b0000000100000110_0;
      patterns[896] = 17'b1000001000000000_0;
      patterns[897] = 17'b1001001000000000_0;
      patterns[898] = 17'b1010001000000000_0;
      patterns[899] = 17'b1011001000000000_0;
      patterns[900] = 17'b0101001000000000_0;
      patterns[901] = 17'b0100001000000000_1;
      patterns[902] = 17'b0000001010101001_0;
      patterns[903] = 17'b1000001000000001_0;
      patterns[904] = 17'b1001001000000001_0;
      patterns[905] = 17'b1010001000000001_0;
      patterns[906] = 17'b1011001000000001_0;
      patterns[907] = 17'b0101001000000000_0;
      patterns[908] = 17'b0100001000000000_1;
      patterns[909] = 17'b0000001000010101_0;
      patterns[910] = 17'b1000001000000010_0;
      patterns[911] = 17'b1001001000000010_0;
      patterns[912] = 17'b1010001000000010_0;
      patterns[913] = 17'b1011001000000010_0;
      patterns[914] = 17'b0101001000000000_0;
      patterns[915] = 17'b0100001000000000_1;
      patterns[916] = 17'b0000001001101011_0;
      patterns[917] = 17'b1000001000000011_0;
      patterns[918] = 17'b1001001000000011_0;
      patterns[919] = 17'b1010001000000011_0;
      patterns[920] = 17'b1011001000000011_0;
      patterns[921] = 17'b0101001000000000_0;
      patterns[922] = 17'b0100001000000000_1;
      patterns[923] = 17'b0000001010001101_0;
      patterns[924] = 17'b1000001000000100_0;
      patterns[925] = 17'b1001001000000100_0;
      patterns[926] = 17'b1010001000000100_0;
      patterns[927] = 17'b1011001000000100_0;
      patterns[928] = 17'b0101001000000000_0;
      patterns[929] = 17'b0100001000000000_1;
      patterns[930] = 17'b0000001001001110_0;
      patterns[931] = 17'b1000001000000101_0;
      patterns[932] = 17'b1001001000000101_0;
      patterns[933] = 17'b1010001000000101_0;
      patterns[934] = 17'b1011001000000101_0;
      patterns[935] = 17'b0101001000000000_0;
      patterns[936] = 17'b0100001000000000_1;
      patterns[937] = 17'b0000001000100111_0;
      patterns[938] = 17'b1000001000000110_0;
      patterns[939] = 17'b1001001000000110_0;
      patterns[940] = 17'b1010001000000110_0;
      patterns[941] = 17'b1011001000000110_0;
      patterns[942] = 17'b0101001000000000_0;
      patterns[943] = 17'b0100001000000000_1;
      patterns[944] = 17'b0000001000111111_0;
      patterns[945] = 17'b1000001000000111_0;
      patterns[946] = 17'b1001001000000111_0;
      patterns[947] = 17'b1010001000000111_0;
      patterns[948] = 17'b1011001000000111_0;
      patterns[949] = 17'b0101001000000000_0;
      patterns[950] = 17'b0100001000000000_1;
      patterns[951] = 17'b0000001011111100_0;
      patterns[952] = 17'b1000001000010000_0;
      patterns[953] = 17'b1001001000010000_0;
      patterns[954] = 17'b1010001000010000_0;
      patterns[955] = 17'b1011001000010000_0;
      patterns[956] = 17'b0101001000010000_0;
      patterns[957] = 17'b0100001000010000_1;
      patterns[958] = 17'b0000001010111100_0;
      patterns[959] = 17'b1000001000010001_0;
      patterns[960] = 17'b1001001000010001_0;
      patterns[961] = 17'b1010001000010001_0;
      patterns[962] = 17'b1011001000010001_0;
      patterns[963] = 17'b0101001000010000_0;
      patterns[964] = 17'b0100001000010000_1;
      patterns[965] = 17'b0000001011101011_0;
      patterns[966] = 17'b1000001000010010_0;
      patterns[967] = 17'b1001001000010010_0;
      patterns[968] = 17'b1010001000010010_0;
      patterns[969] = 17'b1011001000010010_0;
      patterns[970] = 17'b0101001000010000_0;
      patterns[971] = 17'b0100001000010000_1;
      patterns[972] = 17'b0000001001111110_0;
      patterns[973] = 17'b1000001000010011_0;
      patterns[974] = 17'b1001001000010011_0;
      patterns[975] = 17'b1010001000010011_0;
      patterns[976] = 17'b1011001000010011_0;
      patterns[977] = 17'b0101001000010000_0;
      patterns[978] = 17'b0100001000010000_1;
      patterns[979] = 17'b0000001011101010_0;
      patterns[980] = 17'b1000001000010100_0;
      patterns[981] = 17'b1001001000010100_0;
      patterns[982] = 17'b1010001000010100_0;
      patterns[983] = 17'b1011001000010100_0;
      patterns[984] = 17'b0101001000010000_0;
      patterns[985] = 17'b0100001000010000_1;
      patterns[986] = 17'b0000001010100100_0;
      patterns[987] = 17'b1000001000010101_0;
      patterns[988] = 17'b1001001000010101_0;
      patterns[989] = 17'b1010001000010101_0;
      patterns[990] = 17'b1011001000010101_0;
      patterns[991] = 17'b0101001000010000_0;
      patterns[992] = 17'b0100001000010000_1;
      patterns[993] = 17'b0000001011011001_0;
      patterns[994] = 17'b1000001000010110_0;
      patterns[995] = 17'b1001001000010110_0;
      patterns[996] = 17'b1010001000010110_0;
      patterns[997] = 17'b1011001000010110_0;
      patterns[998] = 17'b0101001000010000_0;
      patterns[999] = 17'b0100001000010000_1;
      patterns[1000] = 17'b0000001011111100_0;
      patterns[1001] = 17'b1000001000010111_0;
      patterns[1002] = 17'b1001001000010111_0;
      patterns[1003] = 17'b1010001000010111_0;
      patterns[1004] = 17'b1011001000010111_0;
      patterns[1005] = 17'b0101001000010000_0;
      patterns[1006] = 17'b0100001000010000_1;
      patterns[1007] = 17'b0000001010010100_0;
      patterns[1008] = 17'b1000001000100000_0;
      patterns[1009] = 17'b1001001000100000_0;
      patterns[1010] = 17'b1010001000100000_0;
      patterns[1011] = 17'b1011001000100000_0;
      patterns[1012] = 17'b0101001000100000_0;
      patterns[1013] = 17'b0100001000100000_1;
      patterns[1014] = 17'b0000001011000000_0;
      patterns[1015] = 17'b1000001000100001_0;
      patterns[1016] = 17'b1001001000100001_0;
      patterns[1017] = 17'b1010001000100001_0;
      patterns[1018] = 17'b1011001000100001_0;
      patterns[1019] = 17'b0101001000100000_0;
      patterns[1020] = 17'b0100001000100000_1;
      patterns[1021] = 17'b0000001011101100_0;
      patterns[1022] = 17'b1000001000100010_0;
      patterns[1023] = 17'b1001001000100010_0;
      patterns[1024] = 17'b1010001000100010_0;
      patterns[1025] = 17'b1011001000100010_0;
      patterns[1026] = 17'b0101001000100000_0;
      patterns[1027] = 17'b0100001000100000_1;
      patterns[1028] = 17'b0000001000101101_0;
      patterns[1029] = 17'b1000001000100011_0;
      patterns[1030] = 17'b1001001000100011_0;
      patterns[1031] = 17'b1010001000100011_0;
      patterns[1032] = 17'b1011001000100011_0;
      patterns[1033] = 17'b0101001000100000_0;
      patterns[1034] = 17'b0100001000100000_1;
      patterns[1035] = 17'b0000001001010111_0;
      patterns[1036] = 17'b1000001000100100_0;
      patterns[1037] = 17'b1001001000100100_0;
      patterns[1038] = 17'b1010001000100100_0;
      patterns[1039] = 17'b1011001000100100_0;
      patterns[1040] = 17'b0101001000100000_0;
      patterns[1041] = 17'b0100001000100000_1;
      patterns[1042] = 17'b0000001000111101_0;
      patterns[1043] = 17'b1000001000100101_0;
      patterns[1044] = 17'b1001001000100101_0;
      patterns[1045] = 17'b1010001000100101_0;
      patterns[1046] = 17'b1011001000100101_0;
      patterns[1047] = 17'b0101001000100000_0;
      patterns[1048] = 17'b0100001000100000_1;
      patterns[1049] = 17'b0000001010000011_0;
      patterns[1050] = 17'b1000001000100110_0;
      patterns[1051] = 17'b1001001000100110_0;
      patterns[1052] = 17'b1010001000100110_0;
      patterns[1053] = 17'b1011001000100110_0;
      patterns[1054] = 17'b0101001000100000_0;
      patterns[1055] = 17'b0100001000100000_1;
      patterns[1056] = 17'b0000001011110010_0;
      patterns[1057] = 17'b1000001000100111_0;
      patterns[1058] = 17'b1001001000100111_0;
      patterns[1059] = 17'b1010001000100111_0;
      patterns[1060] = 17'b1011001000100111_0;
      patterns[1061] = 17'b0101001000100000_0;
      patterns[1062] = 17'b0100001000100000_1;
      patterns[1063] = 17'b0000001001000011_0;
      patterns[1064] = 17'b1000001000110000_0;
      patterns[1065] = 17'b1001001000110000_0;
      patterns[1066] = 17'b1010001000110000_0;
      patterns[1067] = 17'b1011001000110000_0;
      patterns[1068] = 17'b0101001000110000_0;
      patterns[1069] = 17'b0100001000110000_1;
      patterns[1070] = 17'b0000001000110010_0;
      patterns[1071] = 17'b1000001000110001_0;
      patterns[1072] = 17'b1001001000110001_0;
      patterns[1073] = 17'b1010001000110001_0;
      patterns[1074] = 17'b1011001000110001_0;
      patterns[1075] = 17'b0101001000110000_0;
      patterns[1076] = 17'b0100001000110000_1;
      patterns[1077] = 17'b0000001001100011_0;
      patterns[1078] = 17'b1000001000110010_0;
      patterns[1079] = 17'b1001001000110010_0;
      patterns[1080] = 17'b1010001000110010_0;
      patterns[1081] = 17'b1011001000110010_0;
      patterns[1082] = 17'b0101001000110000_0;
      patterns[1083] = 17'b0100001000110000_1;
      patterns[1084] = 17'b0000001000000110_0;
      patterns[1085] = 17'b1000001000110011_0;
      patterns[1086] = 17'b1001001000110011_0;
      patterns[1087] = 17'b1010001000110011_0;
      patterns[1088] = 17'b1011001000110011_0;
      patterns[1089] = 17'b0101001000110000_0;
      patterns[1090] = 17'b0100001000110000_1;
      patterns[1091] = 17'b0000001001100110_0;
      patterns[1092] = 17'b1000001000110100_0;
      patterns[1093] = 17'b1001001000110100_0;
      patterns[1094] = 17'b1010001000110100_0;
      patterns[1095] = 17'b1011001000110100_0;
      patterns[1096] = 17'b0101001000110000_0;
      patterns[1097] = 17'b0100001000110000_1;
      patterns[1098] = 17'b0000001000101001_0;
      patterns[1099] = 17'b1000001000110101_0;
      patterns[1100] = 17'b1001001000110101_0;
      patterns[1101] = 17'b1010001000110101_0;
      patterns[1102] = 17'b1011001000110101_0;
      patterns[1103] = 17'b0101001000110000_0;
      patterns[1104] = 17'b0100001000110000_1;
      patterns[1105] = 17'b0000001010111011_0;
      patterns[1106] = 17'b1000001000110110_0;
      patterns[1107] = 17'b1001001000110110_0;
      patterns[1108] = 17'b1010001000110110_0;
      patterns[1109] = 17'b1011001000110110_0;
      patterns[1110] = 17'b0101001000110000_0;
      patterns[1111] = 17'b0100001000110000_1;
      patterns[1112] = 17'b0000001011110101_0;
      patterns[1113] = 17'b1000001000110111_0;
      patterns[1114] = 17'b1001001000110111_0;
      patterns[1115] = 17'b1010001000110111_0;
      patterns[1116] = 17'b1011001000110111_0;
      patterns[1117] = 17'b0101001000110000_0;
      patterns[1118] = 17'b0100001000110000_1;
      patterns[1119] = 17'b0000001010010111_0;
      patterns[1120] = 17'b1000001001000000_0;
      patterns[1121] = 17'b1001001001000000_0;
      patterns[1122] = 17'b1010001001000000_0;
      patterns[1123] = 17'b1011001001000000_0;
      patterns[1124] = 17'b0101001001000000_0;
      patterns[1125] = 17'b0100001001000000_1;
      patterns[1126] = 17'b0000001000101011_0;
      patterns[1127] = 17'b1000001001000001_0;
      patterns[1128] = 17'b1001001001000001_0;
      patterns[1129] = 17'b1010001001000001_0;
      patterns[1130] = 17'b1011001001000001_0;
      patterns[1131] = 17'b0101001001000000_0;
      patterns[1132] = 17'b0100001001000000_1;
      patterns[1133] = 17'b0000001010000011_0;
      patterns[1134] = 17'b1000001001000010_0;
      patterns[1135] = 17'b1001001001000010_0;
      patterns[1136] = 17'b1010001001000010_0;
      patterns[1137] = 17'b1011001001000010_0;
      patterns[1138] = 17'b0101001001000000_0;
      patterns[1139] = 17'b0100001001000000_1;
      patterns[1140] = 17'b0000001001111100_0;
      patterns[1141] = 17'b1000001001000011_0;
      patterns[1142] = 17'b1001001001000011_0;
      patterns[1143] = 17'b1010001001000011_0;
      patterns[1144] = 17'b1011001001000011_0;
      patterns[1145] = 17'b0101001001000000_0;
      patterns[1146] = 17'b0100001001000000_1;
      patterns[1147] = 17'b0000001010101101_0;
      patterns[1148] = 17'b1000001001000100_0;
      patterns[1149] = 17'b1001001001000100_0;
      patterns[1150] = 17'b1010001001000100_0;
      patterns[1151] = 17'b1011001001000100_0;
      patterns[1152] = 17'b0101001001000000_0;
      patterns[1153] = 17'b0100001001000000_1;
      patterns[1154] = 17'b0000001001011010_0;
      patterns[1155] = 17'b1000001001000101_0;
      patterns[1156] = 17'b1001001001000101_0;
      patterns[1157] = 17'b1010001001000101_0;
      patterns[1158] = 17'b1011001001000101_0;
      patterns[1159] = 17'b0101001001000000_0;
      patterns[1160] = 17'b0100001001000000_1;
      patterns[1161] = 17'b0000001000000101_0;
      patterns[1162] = 17'b1000001001000110_0;
      patterns[1163] = 17'b1001001001000110_0;
      patterns[1164] = 17'b1010001001000110_0;
      patterns[1165] = 17'b1011001001000110_0;
      patterns[1166] = 17'b0101001001000000_0;
      patterns[1167] = 17'b0100001001000000_1;
      patterns[1168] = 17'b0000001001011010_0;
      patterns[1169] = 17'b1000001001000111_0;
      patterns[1170] = 17'b1001001001000111_0;
      patterns[1171] = 17'b1010001001000111_0;
      patterns[1172] = 17'b1011001001000111_0;
      patterns[1173] = 17'b0101001001000000_0;
      patterns[1174] = 17'b0100001001000000_1;
      patterns[1175] = 17'b0000001000101011_0;
      patterns[1176] = 17'b1000001001010000_0;
      patterns[1177] = 17'b1001001001010000_0;
      patterns[1178] = 17'b1010001001010000_0;
      patterns[1179] = 17'b1011001001010000_0;
      patterns[1180] = 17'b0101001001010000_0;
      patterns[1181] = 17'b0100001001010000_1;
      patterns[1182] = 17'b0000001001000000_0;
      patterns[1183] = 17'b1000001001010001_0;
      patterns[1184] = 17'b1001001001010001_0;
      patterns[1185] = 17'b1010001001010001_0;
      patterns[1186] = 17'b1011001001010001_0;
      patterns[1187] = 17'b0101001001010000_0;
      patterns[1188] = 17'b0100001001010000_1;
      patterns[1189] = 17'b0000001000010011_0;
      patterns[1190] = 17'b1000001001010010_0;
      patterns[1191] = 17'b1001001001010010_0;
      patterns[1192] = 17'b1010001001010010_0;
      patterns[1193] = 17'b1011001001010010_0;
      patterns[1194] = 17'b0101001001010000_0;
      patterns[1195] = 17'b0100001001010000_1;
      patterns[1196] = 17'b0000001000011101_0;
      patterns[1197] = 17'b1000001001010011_0;
      patterns[1198] = 17'b1001001001010011_0;
      patterns[1199] = 17'b1010001001010011_0;
      patterns[1200] = 17'b1011001001010011_0;
      patterns[1201] = 17'b0101001001010000_0;
      patterns[1202] = 17'b0100001001010000_1;
      patterns[1203] = 17'b0000001011010001_0;
      patterns[1204] = 17'b1000001001010100_0;
      patterns[1205] = 17'b1001001001010100_0;
      patterns[1206] = 17'b1010001001010100_0;
      patterns[1207] = 17'b1011001001010100_0;
      patterns[1208] = 17'b0101001001010000_0;
      patterns[1209] = 17'b0100001001010000_1;
      patterns[1210] = 17'b0000001000001101_0;
      patterns[1211] = 17'b1000001001010101_0;
      patterns[1212] = 17'b1001001001010101_0;
      patterns[1213] = 17'b1010001001010101_0;
      patterns[1214] = 17'b1011001001010101_0;
      patterns[1215] = 17'b0101001001010000_0;
      patterns[1216] = 17'b0100001001010000_1;
      patterns[1217] = 17'b0000001011101111_0;
      patterns[1218] = 17'b1000001001010110_0;
      patterns[1219] = 17'b1001001001010110_0;
      patterns[1220] = 17'b1010001001010110_0;
      patterns[1221] = 17'b1011001001010110_0;
      patterns[1222] = 17'b0101001001010000_0;
      patterns[1223] = 17'b0100001001010000_1;
      patterns[1224] = 17'b0000001000111100_0;
      patterns[1225] = 17'b1000001001010111_0;
      patterns[1226] = 17'b1001001001010111_0;
      patterns[1227] = 17'b1010001001010111_0;
      patterns[1228] = 17'b1011001001010111_0;
      patterns[1229] = 17'b0101001001010000_0;
      patterns[1230] = 17'b0100001001010000_1;
      patterns[1231] = 17'b0000001001101000_0;
      patterns[1232] = 17'b1000001001100000_0;
      patterns[1233] = 17'b1001001001100000_0;
      patterns[1234] = 17'b1010001001100000_0;
      patterns[1235] = 17'b1011001001100000_0;
      patterns[1236] = 17'b0101001001100000_0;
      patterns[1237] = 17'b0100001001100000_1;
      patterns[1238] = 17'b0000001010111010_0;
      patterns[1239] = 17'b1000001001100001_0;
      patterns[1240] = 17'b1001001001100001_0;
      patterns[1241] = 17'b1010001001100001_0;
      patterns[1242] = 17'b1011001001100001_0;
      patterns[1243] = 17'b0101001001100000_0;
      patterns[1244] = 17'b0100001001100000_1;
      patterns[1245] = 17'b0000001010001110_0;
      patterns[1246] = 17'b1000001001100010_0;
      patterns[1247] = 17'b1001001001100010_0;
      patterns[1248] = 17'b1010001001100010_0;
      patterns[1249] = 17'b1011001001100010_0;
      patterns[1250] = 17'b0101001001100000_0;
      patterns[1251] = 17'b0100001001100000_1;
      patterns[1252] = 17'b0000001011010001_0;
      patterns[1253] = 17'b1000001001100011_0;
      patterns[1254] = 17'b1001001001100011_0;
      patterns[1255] = 17'b1010001001100011_0;
      patterns[1256] = 17'b1011001001100011_0;
      patterns[1257] = 17'b0101001001100000_0;
      patterns[1258] = 17'b0100001001100000_1;
      patterns[1259] = 17'b0000001011011100_0;
      patterns[1260] = 17'b1000001001100100_0;
      patterns[1261] = 17'b1001001001100100_0;
      patterns[1262] = 17'b1010001001100100_0;
      patterns[1263] = 17'b1011001001100100_0;
      patterns[1264] = 17'b0101001001100000_0;
      patterns[1265] = 17'b0100001001100000_1;
      patterns[1266] = 17'b0000001010100110_0;
      patterns[1267] = 17'b1000001001100101_0;
      patterns[1268] = 17'b1001001001100101_0;
      patterns[1269] = 17'b1010001001100101_0;
      patterns[1270] = 17'b1011001001100101_0;
      patterns[1271] = 17'b0101001001100000_0;
      patterns[1272] = 17'b0100001001100000_1;
      patterns[1273] = 17'b0000001010011000_0;
      patterns[1274] = 17'b1000001001100110_0;
      patterns[1275] = 17'b1001001001100110_0;
      patterns[1276] = 17'b1010001001100110_0;
      patterns[1277] = 17'b1011001001100110_0;
      patterns[1278] = 17'b0101001001100000_0;
      patterns[1279] = 17'b0100001001100000_1;
      patterns[1280] = 17'b0000001010101111_0;
      patterns[1281] = 17'b1000001001100111_0;
      patterns[1282] = 17'b1001001001100111_0;
      patterns[1283] = 17'b1010001001100111_0;
      patterns[1284] = 17'b1011001001100111_0;
      patterns[1285] = 17'b0101001001100000_0;
      patterns[1286] = 17'b0100001001100000_1;
      patterns[1287] = 17'b0000001010000111_0;
      patterns[1288] = 17'b1000001001110000_0;
      patterns[1289] = 17'b1001001001110000_0;
      patterns[1290] = 17'b1010001001110000_0;
      patterns[1291] = 17'b1011001001110000_0;
      patterns[1292] = 17'b0101001001110000_0;
      patterns[1293] = 17'b0100001001110000_1;
      patterns[1294] = 17'b0000001001111100_0;
      patterns[1295] = 17'b1000001001110001_0;
      patterns[1296] = 17'b1001001001110001_0;
      patterns[1297] = 17'b1010001001110001_0;
      patterns[1298] = 17'b1011001001110001_0;
      patterns[1299] = 17'b0101001001110000_0;
      patterns[1300] = 17'b0100001001110000_1;
      patterns[1301] = 17'b0000001000101111_0;
      patterns[1302] = 17'b1000001001110010_0;
      patterns[1303] = 17'b1001001001110010_0;
      patterns[1304] = 17'b1010001001110010_0;
      patterns[1305] = 17'b1011001001110010_0;
      patterns[1306] = 17'b0101001001110000_0;
      patterns[1307] = 17'b0100001001110000_1;
      patterns[1308] = 17'b0000001000001010_0;
      patterns[1309] = 17'b1000001001110011_0;
      patterns[1310] = 17'b1001001001110011_0;
      patterns[1311] = 17'b1010001001110011_0;
      patterns[1312] = 17'b1011001001110011_0;
      patterns[1313] = 17'b0101001001110000_0;
      patterns[1314] = 17'b0100001001110000_1;
      patterns[1315] = 17'b0000001001010101_0;
      patterns[1316] = 17'b1000001001110100_0;
      patterns[1317] = 17'b1001001001110100_0;
      patterns[1318] = 17'b1010001001110100_0;
      patterns[1319] = 17'b1011001001110100_0;
      patterns[1320] = 17'b0101001001110000_0;
      patterns[1321] = 17'b0100001001110000_1;
      patterns[1322] = 17'b0000001010000110_0;
      patterns[1323] = 17'b1000001001110101_0;
      patterns[1324] = 17'b1001001001110101_0;
      patterns[1325] = 17'b1010001001110101_0;
      patterns[1326] = 17'b1011001001110101_0;
      patterns[1327] = 17'b0101001001110000_0;
      patterns[1328] = 17'b0100001001110000_1;
      patterns[1329] = 17'b0000001000111001_0;
      patterns[1330] = 17'b1000001001110110_0;
      patterns[1331] = 17'b1001001001110110_0;
      patterns[1332] = 17'b1010001001110110_0;
      patterns[1333] = 17'b1011001001110110_0;
      patterns[1334] = 17'b0101001001110000_0;
      patterns[1335] = 17'b0100001001110000_1;
      patterns[1336] = 17'b0000001011110110_0;
      patterns[1337] = 17'b1000001001110111_0;
      patterns[1338] = 17'b1001001001110111_0;
      patterns[1339] = 17'b1010001001110111_0;
      patterns[1340] = 17'b1011001001110111_0;
      patterns[1341] = 17'b0101001001110000_0;
      patterns[1342] = 17'b0100001001110000_1;
      patterns[1343] = 17'b0000001001111001_0;
      patterns[1344] = 17'b1000001100000000_0;
      patterns[1345] = 17'b1001001100000000_0;
      patterns[1346] = 17'b1010001100000000_0;
      patterns[1347] = 17'b1011001100000000_0;
      patterns[1348] = 17'b0101001100000000_0;
      patterns[1349] = 17'b0100001100000000_1;
      patterns[1350] = 17'b0000001100110010_0;
      patterns[1351] = 17'b1000001100000001_0;
      patterns[1352] = 17'b1001001100000001_0;
      patterns[1353] = 17'b1010001100000001_0;
      patterns[1354] = 17'b1011001100000001_0;
      patterns[1355] = 17'b0101001100000000_0;
      patterns[1356] = 17'b0100001100000000_1;
      patterns[1357] = 17'b0000001110111110_0;
      patterns[1358] = 17'b1000001100000010_0;
      patterns[1359] = 17'b1001001100000010_0;
      patterns[1360] = 17'b1010001100000010_0;
      patterns[1361] = 17'b1011001100000010_0;
      patterns[1362] = 17'b0101001100000000_0;
      patterns[1363] = 17'b0100001100000000_1;
      patterns[1364] = 17'b0000001100001001_0;
      patterns[1365] = 17'b1000001100000011_0;
      patterns[1366] = 17'b1001001100000011_0;
      patterns[1367] = 17'b1010001100000011_0;
      patterns[1368] = 17'b1011001100000011_0;
      patterns[1369] = 17'b0101001100000000_0;
      patterns[1370] = 17'b0100001100000000_1;
      patterns[1371] = 17'b0000001111111100_0;
      patterns[1372] = 17'b1000001100000100_0;
      patterns[1373] = 17'b1001001100000100_0;
      patterns[1374] = 17'b1010001100000100_0;
      patterns[1375] = 17'b1011001100000100_0;
      patterns[1376] = 17'b0101001100000000_0;
      patterns[1377] = 17'b0100001100000000_1;
      patterns[1378] = 17'b0000001110001110_0;
      patterns[1379] = 17'b1000001100000101_0;
      patterns[1380] = 17'b1001001100000101_0;
      patterns[1381] = 17'b1010001100000101_0;
      patterns[1382] = 17'b1011001100000101_0;
      patterns[1383] = 17'b0101001100000000_0;
      patterns[1384] = 17'b0100001100000000_1;
      patterns[1385] = 17'b0000001110101001_0;
      patterns[1386] = 17'b1000001100000110_0;
      patterns[1387] = 17'b1001001100000110_0;
      patterns[1388] = 17'b1010001100000110_0;
      patterns[1389] = 17'b1011001100000110_0;
      patterns[1390] = 17'b0101001100000000_0;
      patterns[1391] = 17'b0100001100000000_1;
      patterns[1392] = 17'b0000001111110110_0;
      patterns[1393] = 17'b1000001100000111_0;
      patterns[1394] = 17'b1001001100000111_0;
      patterns[1395] = 17'b1010001100000111_0;
      patterns[1396] = 17'b1011001100000111_0;
      patterns[1397] = 17'b0101001100000000_0;
      patterns[1398] = 17'b0100001100000000_1;
      patterns[1399] = 17'b0000001110111111_0;
      patterns[1400] = 17'b1000001100010000_0;
      patterns[1401] = 17'b1001001100010000_0;
      patterns[1402] = 17'b1010001100010000_0;
      patterns[1403] = 17'b1011001100010000_0;
      patterns[1404] = 17'b0101001100010000_0;
      patterns[1405] = 17'b0100001100010000_1;
      patterns[1406] = 17'b0000001110101000_0;
      patterns[1407] = 17'b1000001100010001_0;
      patterns[1408] = 17'b1001001100010001_0;
      patterns[1409] = 17'b1010001100010001_0;
      patterns[1410] = 17'b1011001100010001_0;
      patterns[1411] = 17'b0101001100010000_0;
      patterns[1412] = 17'b0100001100010000_1;
      patterns[1413] = 17'b0000001100001011_0;
      patterns[1414] = 17'b1000001100010010_0;
      patterns[1415] = 17'b1001001100010010_0;
      patterns[1416] = 17'b1010001100010010_0;
      patterns[1417] = 17'b1011001100010010_0;
      patterns[1418] = 17'b0101001100010000_0;
      patterns[1419] = 17'b0100001100010000_1;
      patterns[1420] = 17'b0000001110101010_0;
      patterns[1421] = 17'b1000001100010011_0;
      patterns[1422] = 17'b1001001100010011_0;
      patterns[1423] = 17'b1010001100010011_0;
      patterns[1424] = 17'b1011001100010011_0;
      patterns[1425] = 17'b0101001100010000_0;
      patterns[1426] = 17'b0100001100010000_1;
      patterns[1427] = 17'b0000001100110110_0;
      patterns[1428] = 17'b1000001100010100_0;
      patterns[1429] = 17'b1001001100010100_0;
      patterns[1430] = 17'b1010001100010100_0;
      patterns[1431] = 17'b1011001100010100_0;
      patterns[1432] = 17'b0101001100010000_0;
      patterns[1433] = 17'b0100001100010000_1;
      patterns[1434] = 17'b0000001101001000_0;
      patterns[1435] = 17'b1000001100010101_0;
      patterns[1436] = 17'b1001001100010101_0;
      patterns[1437] = 17'b1010001100010101_0;
      patterns[1438] = 17'b1011001100010101_0;
      patterns[1439] = 17'b0101001100010000_0;
      patterns[1440] = 17'b0100001100010000_1;
      patterns[1441] = 17'b0000001111100111_0;
      patterns[1442] = 17'b1000001100010110_0;
      patterns[1443] = 17'b1001001100010110_0;
      patterns[1444] = 17'b1010001100010110_0;
      patterns[1445] = 17'b1011001100010110_0;
      patterns[1446] = 17'b0101001100010000_0;
      patterns[1447] = 17'b0100001100010000_1;
      patterns[1448] = 17'b0000001110000000_0;
      patterns[1449] = 17'b1000001100010111_0;
      patterns[1450] = 17'b1001001100010111_0;
      patterns[1451] = 17'b1010001100010111_0;
      patterns[1452] = 17'b1011001100010111_0;
      patterns[1453] = 17'b0101001100010000_0;
      patterns[1454] = 17'b0100001100010000_1;
      patterns[1455] = 17'b0000001100111111_0;
      patterns[1456] = 17'b1000001100100000_0;
      patterns[1457] = 17'b1001001100100000_0;
      patterns[1458] = 17'b1010001100100000_0;
      patterns[1459] = 17'b1011001100100000_0;
      patterns[1460] = 17'b0101001100100000_0;
      patterns[1461] = 17'b0100001100100000_1;
      patterns[1462] = 17'b0000001101010001_0;
      patterns[1463] = 17'b1000001100100001_0;
      patterns[1464] = 17'b1001001100100001_0;
      patterns[1465] = 17'b1010001100100001_0;
      patterns[1466] = 17'b1011001100100001_0;
      patterns[1467] = 17'b0101001100100000_0;
      patterns[1468] = 17'b0100001100100000_1;
      patterns[1469] = 17'b0000001101100000_0;
      patterns[1470] = 17'b1000001100100010_0;
      patterns[1471] = 17'b1001001100100010_0;
      patterns[1472] = 17'b1010001100100010_0;
      patterns[1473] = 17'b1011001100100010_0;
      patterns[1474] = 17'b0101001100100000_0;
      patterns[1475] = 17'b0100001100100000_1;
      patterns[1476] = 17'b0000001101011100_0;
      patterns[1477] = 17'b1000001100100011_0;
      patterns[1478] = 17'b1001001100100011_0;
      patterns[1479] = 17'b1010001100100011_0;
      patterns[1480] = 17'b1011001100100011_0;
      patterns[1481] = 17'b0101001100100000_0;
      patterns[1482] = 17'b0100001100100000_1;
      patterns[1483] = 17'b0000001101111100_0;
      patterns[1484] = 17'b1000001100100100_0;
      patterns[1485] = 17'b1001001100100100_0;
      patterns[1486] = 17'b1010001100100100_0;
      patterns[1487] = 17'b1011001100100100_0;
      patterns[1488] = 17'b0101001100100000_0;
      patterns[1489] = 17'b0100001100100000_1;
      patterns[1490] = 17'b0000001111110000_0;
      patterns[1491] = 17'b1000001100100101_0;
      patterns[1492] = 17'b1001001100100101_0;
      patterns[1493] = 17'b1010001100100101_0;
      patterns[1494] = 17'b1011001100100101_0;
      patterns[1495] = 17'b0101001100100000_0;
      patterns[1496] = 17'b0100001100100000_1;
      patterns[1497] = 17'b0000001100010110_0;
      patterns[1498] = 17'b1000001100100110_0;
      patterns[1499] = 17'b1001001100100110_0;
      patterns[1500] = 17'b1010001100100110_0;
      patterns[1501] = 17'b1011001100100110_0;
      patterns[1502] = 17'b0101001100100000_0;
      patterns[1503] = 17'b0100001100100000_1;
      patterns[1504] = 17'b0000001100110001_0;
      patterns[1505] = 17'b1000001100100111_0;
      patterns[1506] = 17'b1001001100100111_0;
      patterns[1507] = 17'b1010001100100111_0;
      patterns[1508] = 17'b1011001100100111_0;
      patterns[1509] = 17'b0101001100100000_0;
      patterns[1510] = 17'b0100001100100000_1;
      patterns[1511] = 17'b0000001110100110_0;
      patterns[1512] = 17'b1000001100110000_0;
      patterns[1513] = 17'b1001001100110000_0;
      patterns[1514] = 17'b1010001100110000_0;
      patterns[1515] = 17'b1011001100110000_0;
      patterns[1516] = 17'b0101001100110000_0;
      patterns[1517] = 17'b0100001100110000_1;
      patterns[1518] = 17'b0000001101110010_0;
      patterns[1519] = 17'b1000001100110001_0;
      patterns[1520] = 17'b1001001100110001_0;
      patterns[1521] = 17'b1010001100110001_0;
      patterns[1522] = 17'b1011001100110001_0;
      patterns[1523] = 17'b0101001100110000_0;
      patterns[1524] = 17'b0100001100110000_1;
      patterns[1525] = 17'b0000001101101110_0;
      patterns[1526] = 17'b1000001100110010_0;
      patterns[1527] = 17'b1001001100110010_0;
      patterns[1528] = 17'b1010001100110010_0;
      patterns[1529] = 17'b1011001100110010_0;
      patterns[1530] = 17'b0101001100110000_0;
      patterns[1531] = 17'b0100001100110000_1;
      patterns[1532] = 17'b0000001100101001_0;
      patterns[1533] = 17'b1000001100110011_0;
      patterns[1534] = 17'b1001001100110011_0;
      patterns[1535] = 17'b1010001100110011_0;
      patterns[1536] = 17'b1011001100110011_0;
      patterns[1537] = 17'b0101001100110000_0;
      patterns[1538] = 17'b0100001100110000_1;
      patterns[1539] = 17'b0000001101010111_0;
      patterns[1540] = 17'b1000001100110100_0;
      patterns[1541] = 17'b1001001100110100_0;
      patterns[1542] = 17'b1010001100110100_0;
      patterns[1543] = 17'b1011001100110100_0;
      patterns[1544] = 17'b0101001100110000_0;
      patterns[1545] = 17'b0100001100110000_1;
      patterns[1546] = 17'b0000001111010100_0;
      patterns[1547] = 17'b1000001100110101_0;
      patterns[1548] = 17'b1001001100110101_0;
      patterns[1549] = 17'b1010001100110101_0;
      patterns[1550] = 17'b1011001100110101_0;
      patterns[1551] = 17'b0101001100110000_0;
      patterns[1552] = 17'b0100001100110000_1;
      patterns[1553] = 17'b0000001110000101_0;
      patterns[1554] = 17'b1000001100110110_0;
      patterns[1555] = 17'b1001001100110110_0;
      patterns[1556] = 17'b1010001100110110_0;
      patterns[1557] = 17'b1011001100110110_0;
      patterns[1558] = 17'b0101001100110000_0;
      patterns[1559] = 17'b0100001100110000_1;
      patterns[1560] = 17'b0000001111110001_0;
      patterns[1561] = 17'b1000001100110111_0;
      patterns[1562] = 17'b1001001100110111_0;
      patterns[1563] = 17'b1010001100110111_0;
      patterns[1564] = 17'b1011001100110111_0;
      patterns[1565] = 17'b0101001100110000_0;
      patterns[1566] = 17'b0100001100110000_1;
      patterns[1567] = 17'b0000001100000000_0;
      patterns[1568] = 17'b1000001101000000_0;
      patterns[1569] = 17'b1001001101000000_0;
      patterns[1570] = 17'b1010001101000000_0;
      patterns[1571] = 17'b1011001101000000_0;
      patterns[1572] = 17'b0101001101000000_0;
      patterns[1573] = 17'b0100001101000000_1;
      patterns[1574] = 17'b0000001101101001_0;
      patterns[1575] = 17'b1000001101000001_0;
      patterns[1576] = 17'b1001001101000001_0;
      patterns[1577] = 17'b1010001101000001_0;
      patterns[1578] = 17'b1011001101000001_0;
      patterns[1579] = 17'b0101001101000000_0;
      patterns[1580] = 17'b0100001101000000_1;
      patterns[1581] = 17'b0000001101110001_0;
      patterns[1582] = 17'b1000001101000010_0;
      patterns[1583] = 17'b1001001101000010_0;
      patterns[1584] = 17'b1010001101000010_0;
      patterns[1585] = 17'b1011001101000010_0;
      patterns[1586] = 17'b0101001101000000_0;
      patterns[1587] = 17'b0100001101000000_1;
      patterns[1588] = 17'b0000001111111111_0;
      patterns[1589] = 17'b1000001101000011_0;
      patterns[1590] = 17'b1001001101000011_0;
      patterns[1591] = 17'b1010001101000011_0;
      patterns[1592] = 17'b1011001101000011_0;
      patterns[1593] = 17'b0101001101000000_0;
      patterns[1594] = 17'b0100001101000000_1;
      patterns[1595] = 17'b0000001111000111_0;
      patterns[1596] = 17'b1000001101000100_0;
      patterns[1597] = 17'b1001001101000100_0;
      patterns[1598] = 17'b1010001101000100_0;
      patterns[1599] = 17'b1011001101000100_0;
      patterns[1600] = 17'b0101001101000000_0;
      patterns[1601] = 17'b0100001101000000_1;
      patterns[1602] = 17'b0000001111001010_0;
      patterns[1603] = 17'b1000001101000101_0;
      patterns[1604] = 17'b1001001101000101_0;
      patterns[1605] = 17'b1010001101000101_0;
      patterns[1606] = 17'b1011001101000101_0;
      patterns[1607] = 17'b0101001101000000_0;
      patterns[1608] = 17'b0100001101000000_1;
      patterns[1609] = 17'b0000001110110011_0;
      patterns[1610] = 17'b1000001101000110_0;
      patterns[1611] = 17'b1001001101000110_0;
      patterns[1612] = 17'b1010001101000110_0;
      patterns[1613] = 17'b1011001101000110_0;
      patterns[1614] = 17'b0101001101000000_0;
      patterns[1615] = 17'b0100001101000000_1;
      patterns[1616] = 17'b0000001101011110_0;
      patterns[1617] = 17'b1000001101000111_0;
      patterns[1618] = 17'b1001001101000111_0;
      patterns[1619] = 17'b1010001101000111_0;
      patterns[1620] = 17'b1011001101000111_0;
      patterns[1621] = 17'b0101001101000000_0;
      patterns[1622] = 17'b0100001101000000_1;
      patterns[1623] = 17'b0000001101100110_0;
      patterns[1624] = 17'b1000001101010000_0;
      patterns[1625] = 17'b1001001101010000_0;
      patterns[1626] = 17'b1010001101010000_0;
      patterns[1627] = 17'b1011001101010000_0;
      patterns[1628] = 17'b0101001101010000_0;
      patterns[1629] = 17'b0100001101010000_1;
      patterns[1630] = 17'b0000001100001010_0;
      patterns[1631] = 17'b1000001101010001_0;
      patterns[1632] = 17'b1001001101010001_0;
      patterns[1633] = 17'b1010001101010001_0;
      patterns[1634] = 17'b1011001101010001_0;
      patterns[1635] = 17'b0101001101010000_0;
      patterns[1636] = 17'b0100001101010000_1;
      patterns[1637] = 17'b0000001110001111_0;
      patterns[1638] = 17'b1000001101010010_0;
      patterns[1639] = 17'b1001001101010010_0;
      patterns[1640] = 17'b1010001101010010_0;
      patterns[1641] = 17'b1011001101010010_0;
      patterns[1642] = 17'b0101001101010000_0;
      patterns[1643] = 17'b0100001101010000_1;
      patterns[1644] = 17'b0000001110011111_0;
      patterns[1645] = 17'b1000001101010011_0;
      patterns[1646] = 17'b1001001101010011_0;
      patterns[1647] = 17'b1010001101010011_0;
      patterns[1648] = 17'b1011001101010011_0;
      patterns[1649] = 17'b0101001101010000_0;
      patterns[1650] = 17'b0100001101010000_1;
      patterns[1651] = 17'b0000001100010100_0;
      patterns[1652] = 17'b1000001101010100_0;
      patterns[1653] = 17'b1001001101010100_0;
      patterns[1654] = 17'b1010001101010100_0;
      patterns[1655] = 17'b1011001101010100_0;
      patterns[1656] = 17'b0101001101010000_0;
      patterns[1657] = 17'b0100001101010000_1;
      patterns[1658] = 17'b0000001110101011_0;
      patterns[1659] = 17'b1000001101010101_0;
      patterns[1660] = 17'b1001001101010101_0;
      patterns[1661] = 17'b1010001101010101_0;
      patterns[1662] = 17'b1011001101010101_0;
      patterns[1663] = 17'b0101001101010000_0;
      patterns[1664] = 17'b0100001101010000_1;
      patterns[1665] = 17'b0000001101011001_0;
      patterns[1666] = 17'b1000001101010110_0;
      patterns[1667] = 17'b1001001101010110_0;
      patterns[1668] = 17'b1010001101010110_0;
      patterns[1669] = 17'b1011001101010110_0;
      patterns[1670] = 17'b0101001101010000_0;
      patterns[1671] = 17'b0100001101010000_1;
      patterns[1672] = 17'b0000001110101001_0;
      patterns[1673] = 17'b1000001101010111_0;
      patterns[1674] = 17'b1001001101010111_0;
      patterns[1675] = 17'b1010001101010111_0;
      patterns[1676] = 17'b1011001101010111_0;
      patterns[1677] = 17'b0101001101010000_0;
      patterns[1678] = 17'b0100001101010000_1;
      patterns[1679] = 17'b0000001100010000_0;
      patterns[1680] = 17'b1000001101100000_0;
      patterns[1681] = 17'b1001001101100000_0;
      patterns[1682] = 17'b1010001101100000_0;
      patterns[1683] = 17'b1011001101100000_0;
      patterns[1684] = 17'b0101001101100000_0;
      patterns[1685] = 17'b0100001101100000_1;
      patterns[1686] = 17'b0000001100001100_0;
      patterns[1687] = 17'b1000001101100001_0;
      patterns[1688] = 17'b1001001101100001_0;
      patterns[1689] = 17'b1010001101100001_0;
      patterns[1690] = 17'b1011001101100001_0;
      patterns[1691] = 17'b0101001101100000_0;
      patterns[1692] = 17'b0100001101100000_1;
      patterns[1693] = 17'b0000001110101111_0;
      patterns[1694] = 17'b1000001101100010_0;
      patterns[1695] = 17'b1001001101100010_0;
      patterns[1696] = 17'b1010001101100010_0;
      patterns[1697] = 17'b1011001101100010_0;
      patterns[1698] = 17'b0101001101100000_0;
      patterns[1699] = 17'b0100001101100000_1;
      patterns[1700] = 17'b0000001111011100_0;
      patterns[1701] = 17'b1000001101100011_0;
      patterns[1702] = 17'b1001001101100011_0;
      patterns[1703] = 17'b1010001101100011_0;
      patterns[1704] = 17'b1011001101100011_0;
      patterns[1705] = 17'b0101001101100000_0;
      patterns[1706] = 17'b0100001101100000_1;
      patterns[1707] = 17'b0000001101101011_0;
      patterns[1708] = 17'b1000001101100100_0;
      patterns[1709] = 17'b1001001101100100_0;
      patterns[1710] = 17'b1010001101100100_0;
      patterns[1711] = 17'b1011001101100100_0;
      patterns[1712] = 17'b0101001101100000_0;
      patterns[1713] = 17'b0100001101100000_1;
      patterns[1714] = 17'b0000001100011010_0;
      patterns[1715] = 17'b1000001101100101_0;
      patterns[1716] = 17'b1001001101100101_0;
      patterns[1717] = 17'b1010001101100101_0;
      patterns[1718] = 17'b1011001101100101_0;
      patterns[1719] = 17'b0101001101100000_0;
      patterns[1720] = 17'b0100001101100000_1;
      patterns[1721] = 17'b0000001111110000_0;
      patterns[1722] = 17'b1000001101100110_0;
      patterns[1723] = 17'b1001001101100110_0;
      patterns[1724] = 17'b1010001101100110_0;
      patterns[1725] = 17'b1011001101100110_0;
      patterns[1726] = 17'b0101001101100000_0;
      patterns[1727] = 17'b0100001101100000_1;
      patterns[1728] = 17'b0000001110101110_0;
      patterns[1729] = 17'b1000001101100111_0;
      patterns[1730] = 17'b1001001101100111_0;
      patterns[1731] = 17'b1010001101100111_0;
      patterns[1732] = 17'b1011001101100111_0;
      patterns[1733] = 17'b0101001101100000_0;
      patterns[1734] = 17'b0100001101100000_1;
      patterns[1735] = 17'b0000001100100010_0;
      patterns[1736] = 17'b1000001101110000_0;
      patterns[1737] = 17'b1001001101110000_0;
      patterns[1738] = 17'b1010001101110000_0;
      patterns[1739] = 17'b1011001101110000_0;
      patterns[1740] = 17'b0101001101110000_0;
      patterns[1741] = 17'b0100001101110000_1;
      patterns[1742] = 17'b0000001111111110_0;
      patterns[1743] = 17'b1000001101110001_0;
      patterns[1744] = 17'b1001001101110001_0;
      patterns[1745] = 17'b1010001101110001_0;
      patterns[1746] = 17'b1011001101110001_0;
      patterns[1747] = 17'b0101001101110000_0;
      patterns[1748] = 17'b0100001101110000_1;
      patterns[1749] = 17'b0000001101010010_0;
      patterns[1750] = 17'b1000001101110010_0;
      patterns[1751] = 17'b1001001101110010_0;
      patterns[1752] = 17'b1010001101110010_0;
      patterns[1753] = 17'b1011001101110010_0;
      patterns[1754] = 17'b0101001101110000_0;
      patterns[1755] = 17'b0100001101110000_1;
      patterns[1756] = 17'b0000001100010001_0;
      patterns[1757] = 17'b1000001101110011_0;
      patterns[1758] = 17'b1001001101110011_0;
      patterns[1759] = 17'b1010001101110011_0;
      patterns[1760] = 17'b1011001101110011_0;
      patterns[1761] = 17'b0101001101110000_0;
      patterns[1762] = 17'b0100001101110000_1;
      patterns[1763] = 17'b0000001111010101_0;
      patterns[1764] = 17'b1000001101110100_0;
      patterns[1765] = 17'b1001001101110100_0;
      patterns[1766] = 17'b1010001101110100_0;
      patterns[1767] = 17'b1011001101110100_0;
      patterns[1768] = 17'b0101001101110000_0;
      patterns[1769] = 17'b0100001101110000_1;
      patterns[1770] = 17'b0000001111111110_0;
      patterns[1771] = 17'b1000001101110101_0;
      patterns[1772] = 17'b1001001101110101_0;
      patterns[1773] = 17'b1010001101110101_0;
      patterns[1774] = 17'b1011001101110101_0;
      patterns[1775] = 17'b0101001101110000_0;
      patterns[1776] = 17'b0100001101110000_1;
      patterns[1777] = 17'b0000001101001000_0;
      patterns[1778] = 17'b1000001101110110_0;
      patterns[1779] = 17'b1001001101110110_0;
      patterns[1780] = 17'b1010001101110110_0;
      patterns[1781] = 17'b1011001101110110_0;
      patterns[1782] = 17'b0101001101110000_0;
      patterns[1783] = 17'b0100001101110000_1;
      patterns[1784] = 17'b0000001101010110_0;
      patterns[1785] = 17'b1000001101110111_0;
      patterns[1786] = 17'b1001001101110111_0;
      patterns[1787] = 17'b1010001101110111_0;
      patterns[1788] = 17'b1011001101110111_0;
      patterns[1789] = 17'b0101001101110000_0;
      patterns[1790] = 17'b0100001101110000_1;
      patterns[1791] = 17'b0000001111110010_0;
      patterns[1792] = 17'b1000010000000000_0;
      patterns[1793] = 17'b1001010000000000_0;
      patterns[1794] = 17'b1010010000000000_0;
      patterns[1795] = 17'b1011010000000000_0;
      patterns[1796] = 17'b0101010000000000_0;
      patterns[1797] = 17'b0100010000000000_1;
      patterns[1798] = 17'b0000010001000011_0;
      patterns[1799] = 17'b1000010000000001_0;
      patterns[1800] = 17'b1001010000000001_0;
      patterns[1801] = 17'b1010010000000001_0;
      patterns[1802] = 17'b1011010000000001_0;
      patterns[1803] = 17'b0101010000000000_0;
      patterns[1804] = 17'b0100010000000000_1;
      patterns[1805] = 17'b0000010000100001_0;
      patterns[1806] = 17'b1000010000000010_0;
      patterns[1807] = 17'b1001010000000010_0;
      patterns[1808] = 17'b1010010000000010_0;
      patterns[1809] = 17'b1011010000000010_0;
      patterns[1810] = 17'b0101010000000000_0;
      patterns[1811] = 17'b0100010000000000_1;
      patterns[1812] = 17'b0000010011110110_0;
      patterns[1813] = 17'b1000010000000011_0;
      patterns[1814] = 17'b1001010000000011_0;
      patterns[1815] = 17'b1010010000000011_0;
      patterns[1816] = 17'b1011010000000011_0;
      patterns[1817] = 17'b0101010000000000_0;
      patterns[1818] = 17'b0100010000000000_1;
      patterns[1819] = 17'b0000010001001000_0;
      patterns[1820] = 17'b1000010000000100_0;
      patterns[1821] = 17'b1001010000000100_0;
      patterns[1822] = 17'b1010010000000100_0;
      patterns[1823] = 17'b1011010000000100_0;
      patterns[1824] = 17'b0101010000000000_0;
      patterns[1825] = 17'b0100010000000000_1;
      patterns[1826] = 17'b0000010001110111_0;
      patterns[1827] = 17'b1000010000000101_0;
      patterns[1828] = 17'b1001010000000101_0;
      patterns[1829] = 17'b1010010000000101_0;
      patterns[1830] = 17'b1011010000000101_0;
      patterns[1831] = 17'b0101010000000000_0;
      patterns[1832] = 17'b0100010000000000_1;
      patterns[1833] = 17'b0000010000010011_0;
      patterns[1834] = 17'b1000010000000110_0;
      patterns[1835] = 17'b1001010000000110_0;
      patterns[1836] = 17'b1010010000000110_0;
      patterns[1837] = 17'b1011010000000110_0;
      patterns[1838] = 17'b0101010000000000_0;
      patterns[1839] = 17'b0100010000000000_1;
      patterns[1840] = 17'b0000010010000000_0;
      patterns[1841] = 17'b1000010000000111_0;
      patterns[1842] = 17'b1001010000000111_0;
      patterns[1843] = 17'b1010010000000111_0;
      patterns[1844] = 17'b1011010000000111_0;
      patterns[1845] = 17'b0101010000000000_0;
      patterns[1846] = 17'b0100010000000000_1;
      patterns[1847] = 17'b0000010010111100_0;
      patterns[1848] = 17'b1000010000010000_0;
      patterns[1849] = 17'b1001010000010000_0;
      patterns[1850] = 17'b1010010000010000_0;
      patterns[1851] = 17'b1011010000010000_0;
      patterns[1852] = 17'b0101010000010000_0;
      patterns[1853] = 17'b0100010000010000_1;
      patterns[1854] = 17'b0000010011110111_0;
      patterns[1855] = 17'b1000010000010001_0;
      patterns[1856] = 17'b1001010000010001_0;
      patterns[1857] = 17'b1010010000010001_0;
      patterns[1858] = 17'b1011010000010001_0;
      patterns[1859] = 17'b0101010000010000_0;
      patterns[1860] = 17'b0100010000010000_1;
      patterns[1861] = 17'b0000010000111111_0;
      patterns[1862] = 17'b1000010000010010_0;
      patterns[1863] = 17'b1001010000010010_0;
      patterns[1864] = 17'b1010010000010010_0;
      patterns[1865] = 17'b1011010000010010_0;
      patterns[1866] = 17'b0101010000010000_0;
      patterns[1867] = 17'b0100010000010000_1;
      patterns[1868] = 17'b0000010001001011_0;
      patterns[1869] = 17'b1000010000010011_0;
      patterns[1870] = 17'b1001010000010011_0;
      patterns[1871] = 17'b1010010000010011_0;
      patterns[1872] = 17'b1011010000010011_0;
      patterns[1873] = 17'b0101010000010000_0;
      patterns[1874] = 17'b0100010000010000_1;
      patterns[1875] = 17'b0000010011111110_0;
      patterns[1876] = 17'b1000010000010100_0;
      patterns[1877] = 17'b1001010000010100_0;
      patterns[1878] = 17'b1010010000010100_0;
      patterns[1879] = 17'b1011010000010100_0;
      patterns[1880] = 17'b0101010000010000_0;
      patterns[1881] = 17'b0100010000010000_1;
      patterns[1882] = 17'b0000010001000110_0;
      patterns[1883] = 17'b1000010000010101_0;
      patterns[1884] = 17'b1001010000010101_0;
      patterns[1885] = 17'b1010010000010101_0;
      patterns[1886] = 17'b1011010000010101_0;
      patterns[1887] = 17'b0101010000010000_0;
      patterns[1888] = 17'b0100010000010000_1;
      patterns[1889] = 17'b0000010010001010_0;
      patterns[1890] = 17'b1000010000010110_0;
      patterns[1891] = 17'b1001010000010110_0;
      patterns[1892] = 17'b1010010000010110_0;
      patterns[1893] = 17'b1011010000010110_0;
      patterns[1894] = 17'b0101010000010000_0;
      patterns[1895] = 17'b0100010000010000_1;
      patterns[1896] = 17'b0000010000000100_0;
      patterns[1897] = 17'b1000010000010111_0;
      patterns[1898] = 17'b1001010000010111_0;
      patterns[1899] = 17'b1010010000010111_0;
      patterns[1900] = 17'b1011010000010111_0;
      patterns[1901] = 17'b0101010000010000_0;
      patterns[1902] = 17'b0100010000010000_1;
      patterns[1903] = 17'b0000010011100011_0;
      patterns[1904] = 17'b1000010000100000_0;
      patterns[1905] = 17'b1001010000100000_0;
      patterns[1906] = 17'b1010010000100000_0;
      patterns[1907] = 17'b1011010000100000_0;
      patterns[1908] = 17'b0101010000100000_0;
      patterns[1909] = 17'b0100010000100000_1;
      patterns[1910] = 17'b0000010011011111_0;
      patterns[1911] = 17'b1000010000100001_0;
      patterns[1912] = 17'b1001010000100001_0;
      patterns[1913] = 17'b1010010000100001_0;
      patterns[1914] = 17'b1011010000100001_0;
      patterns[1915] = 17'b0101010000100000_0;
      patterns[1916] = 17'b0100010000100000_1;
      patterns[1917] = 17'b0000010010011000_0;
      patterns[1918] = 17'b1000010000100010_0;
      patterns[1919] = 17'b1001010000100010_0;
      patterns[1920] = 17'b1010010000100010_0;
      patterns[1921] = 17'b1011010000100010_0;
      patterns[1922] = 17'b0101010000100000_0;
      patterns[1923] = 17'b0100010000100000_1;
      patterns[1924] = 17'b0000010011100101_0;
      patterns[1925] = 17'b1000010000100011_0;
      patterns[1926] = 17'b1001010000100011_0;
      patterns[1927] = 17'b1010010000100011_0;
      patterns[1928] = 17'b1011010000100011_0;
      patterns[1929] = 17'b0101010000100000_0;
      patterns[1930] = 17'b0100010000100000_1;
      patterns[1931] = 17'b0000010001001011_0;
      patterns[1932] = 17'b1000010000100100_0;
      patterns[1933] = 17'b1001010000100100_0;
      patterns[1934] = 17'b1010010000100100_0;
      patterns[1935] = 17'b1011010000100100_0;
      patterns[1936] = 17'b0101010000100000_0;
      patterns[1937] = 17'b0100010000100000_1;
      patterns[1938] = 17'b0000010011010010_0;
      patterns[1939] = 17'b1000010000100101_0;
      patterns[1940] = 17'b1001010000100101_0;
      patterns[1941] = 17'b1010010000100101_0;
      patterns[1942] = 17'b1011010000100101_0;
      patterns[1943] = 17'b0101010000100000_0;
      patterns[1944] = 17'b0100010000100000_1;
      patterns[1945] = 17'b0000010010001001_0;
      patterns[1946] = 17'b1000010000100110_0;
      patterns[1947] = 17'b1001010000100110_0;
      patterns[1948] = 17'b1010010000100110_0;
      patterns[1949] = 17'b1011010000100110_0;
      patterns[1950] = 17'b0101010000100000_0;
      patterns[1951] = 17'b0100010000100000_1;
      patterns[1952] = 17'b0000010010011010_0;
      patterns[1953] = 17'b1000010000100111_0;
      patterns[1954] = 17'b1001010000100111_0;
      patterns[1955] = 17'b1010010000100111_0;
      patterns[1956] = 17'b1011010000100111_0;
      patterns[1957] = 17'b0101010000100000_0;
      patterns[1958] = 17'b0100010000100000_1;
      patterns[1959] = 17'b0000010001000111_0;
      patterns[1960] = 17'b1000010000110000_0;
      patterns[1961] = 17'b1001010000110000_0;
      patterns[1962] = 17'b1010010000110000_0;
      patterns[1963] = 17'b1011010000110000_0;
      patterns[1964] = 17'b0101010000110000_0;
      patterns[1965] = 17'b0100010000110000_1;
      patterns[1966] = 17'b0000010010110011_0;
      patterns[1967] = 17'b1000010000110001_0;
      patterns[1968] = 17'b1001010000110001_0;
      patterns[1969] = 17'b1010010000110001_0;
      patterns[1970] = 17'b1011010000110001_0;
      patterns[1971] = 17'b0101010000110000_0;
      patterns[1972] = 17'b0100010000110000_1;
      patterns[1973] = 17'b0000010010101111_0;
      patterns[1974] = 17'b1000010000110010_0;
      patterns[1975] = 17'b1001010000110010_0;
      patterns[1976] = 17'b1010010000110010_0;
      patterns[1977] = 17'b1011010000110010_0;
      patterns[1978] = 17'b0101010000110000_0;
      patterns[1979] = 17'b0100010000110000_1;
      patterns[1980] = 17'b0000010000100101_0;
      patterns[1981] = 17'b1000010000110011_0;
      patterns[1982] = 17'b1001010000110011_0;
      patterns[1983] = 17'b1010010000110011_0;
      patterns[1984] = 17'b1011010000110011_0;
      patterns[1985] = 17'b0101010000110000_0;
      patterns[1986] = 17'b0100010000110000_1;
      patterns[1987] = 17'b0000010010010100_0;
      patterns[1988] = 17'b1000010000110100_0;
      patterns[1989] = 17'b1001010000110100_0;
      patterns[1990] = 17'b1010010000110100_0;
      patterns[1991] = 17'b1011010000110100_0;
      patterns[1992] = 17'b0101010000110000_0;
      patterns[1993] = 17'b0100010000110000_1;
      patterns[1994] = 17'b0000010001010110_0;
      patterns[1995] = 17'b1000010000110101_0;
      patterns[1996] = 17'b1001010000110101_0;
      patterns[1997] = 17'b1010010000110101_0;
      patterns[1998] = 17'b1011010000110101_0;
      patterns[1999] = 17'b0101010000110000_0;
      patterns[2000] = 17'b0100010000110000_1;
      patterns[2001] = 17'b0000010010111110_0;
      patterns[2002] = 17'b1000010000110110_0;
      patterns[2003] = 17'b1001010000110110_0;
      patterns[2004] = 17'b1010010000110110_0;
      patterns[2005] = 17'b1011010000110110_0;
      patterns[2006] = 17'b0101010000110000_0;
      patterns[2007] = 17'b0100010000110000_1;
      patterns[2008] = 17'b0000010010100101_0;
      patterns[2009] = 17'b1000010000110111_0;
      patterns[2010] = 17'b1001010000110111_0;
      patterns[2011] = 17'b1010010000110111_0;
      patterns[2012] = 17'b1011010000110111_0;
      patterns[2013] = 17'b0101010000110000_0;
      patterns[2014] = 17'b0100010000110000_1;
      patterns[2015] = 17'b0000010001001101_0;
      patterns[2016] = 17'b1000010001000000_0;
      patterns[2017] = 17'b1001010001000000_0;
      patterns[2018] = 17'b1010010001000000_0;
      patterns[2019] = 17'b1011010001000000_0;
      patterns[2020] = 17'b0101010001000000_0;
      patterns[2021] = 17'b0100010001000000_1;
      patterns[2022] = 17'b0000010001010101_0;
      patterns[2023] = 17'b1000010001000001_0;
      patterns[2024] = 17'b1001010001000001_0;
      patterns[2025] = 17'b1010010001000001_0;
      patterns[2026] = 17'b1011010001000001_0;
      patterns[2027] = 17'b0101010001000000_0;
      patterns[2028] = 17'b0100010001000000_1;
      patterns[2029] = 17'b0000010010101100_0;
      patterns[2030] = 17'b1000010001000010_0;
      patterns[2031] = 17'b1001010001000010_0;
      patterns[2032] = 17'b1010010001000010_0;
      patterns[2033] = 17'b1011010001000010_0;
      patterns[2034] = 17'b0101010001000000_0;
      patterns[2035] = 17'b0100010001000000_1;
      patterns[2036] = 17'b0000010011110100_0;
      patterns[2037] = 17'b1000010001000011_0;
      patterns[2038] = 17'b1001010001000011_0;
      patterns[2039] = 17'b1010010001000011_0;
      patterns[2040] = 17'b1011010001000011_0;
      patterns[2041] = 17'b0101010001000000_0;
      patterns[2042] = 17'b0100010001000000_1;
      patterns[2043] = 17'b0000010000101110_0;
      patterns[2044] = 17'b1000010001000100_0;
      patterns[2045] = 17'b1001010001000100_0;
      patterns[2046] = 17'b1010010001000100_0;
      patterns[2047] = 17'b1011010001000100_0;
      patterns[2048] = 17'b0101010001000000_0;
      patterns[2049] = 17'b0100010001000000_1;
      patterns[2050] = 17'b0000010011101010_0;
      patterns[2051] = 17'b1000010001000101_0;
      patterns[2052] = 17'b1001010001000101_0;
      patterns[2053] = 17'b1010010001000101_0;
      patterns[2054] = 17'b1011010001000101_0;
      patterns[2055] = 17'b0101010001000000_0;
      patterns[2056] = 17'b0100010001000000_1;
      patterns[2057] = 17'b0000010011011000_0;
      patterns[2058] = 17'b1000010001000110_0;
      patterns[2059] = 17'b1001010001000110_0;
      patterns[2060] = 17'b1010010001000110_0;
      patterns[2061] = 17'b1011010001000110_0;
      patterns[2062] = 17'b0101010001000000_0;
      patterns[2063] = 17'b0100010001000000_1;
      patterns[2064] = 17'b0000010000101101_0;
      patterns[2065] = 17'b1000010001000111_0;
      patterns[2066] = 17'b1001010001000111_0;
      patterns[2067] = 17'b1010010001000111_0;
      patterns[2068] = 17'b1011010001000111_0;
      patterns[2069] = 17'b0101010001000000_0;
      patterns[2070] = 17'b0100010001000000_1;
      patterns[2071] = 17'b0000010010011100_0;
      patterns[2072] = 17'b1000010001010000_0;
      patterns[2073] = 17'b1001010001010000_0;
      patterns[2074] = 17'b1010010001010000_0;
      patterns[2075] = 17'b1011010001010000_0;
      patterns[2076] = 17'b0101010001010000_0;
      patterns[2077] = 17'b0100010001010000_1;
      patterns[2078] = 17'b0000010011100100_0;
      patterns[2079] = 17'b1000010001010001_0;
      patterns[2080] = 17'b1001010001010001_0;
      patterns[2081] = 17'b1010010001010001_0;
      patterns[2082] = 17'b1011010001010001_0;
      patterns[2083] = 17'b0101010001010000_0;
      patterns[2084] = 17'b0100010001010000_1;
      patterns[2085] = 17'b0000010010110011_0;
      patterns[2086] = 17'b1000010001010010_0;
      patterns[2087] = 17'b1001010001010010_0;
      patterns[2088] = 17'b1010010001010010_0;
      patterns[2089] = 17'b1011010001010010_0;
      patterns[2090] = 17'b0101010001010000_0;
      patterns[2091] = 17'b0100010001010000_1;
      patterns[2092] = 17'b0000010010100010_0;
      patterns[2093] = 17'b1000010001010011_0;
      patterns[2094] = 17'b1001010001010011_0;
      patterns[2095] = 17'b1010010001010011_0;
      patterns[2096] = 17'b1011010001010011_0;
      patterns[2097] = 17'b0101010001010000_0;
      patterns[2098] = 17'b0100010001010000_1;
      patterns[2099] = 17'b0000010000111001_0;
      patterns[2100] = 17'b1000010001010100_0;
      patterns[2101] = 17'b1001010001010100_0;
      patterns[2102] = 17'b1010010001010100_0;
      patterns[2103] = 17'b1011010001010100_0;
      patterns[2104] = 17'b0101010001010000_0;
      patterns[2105] = 17'b0100010001010000_1;
      patterns[2106] = 17'b0000010001010110_0;
      patterns[2107] = 17'b1000010001010101_0;
      patterns[2108] = 17'b1001010001010101_0;
      patterns[2109] = 17'b1010010001010101_0;
      patterns[2110] = 17'b1011010001010101_0;
      patterns[2111] = 17'b0101010001010000_0;
      patterns[2112] = 17'b0100010001010000_1;
      patterns[2113] = 17'b0000010011001110_0;
      patterns[2114] = 17'b1000010001010110_0;
      patterns[2115] = 17'b1001010001010110_0;
      patterns[2116] = 17'b1010010001010110_0;
      patterns[2117] = 17'b1011010001010110_0;
      patterns[2118] = 17'b0101010001010000_0;
      patterns[2119] = 17'b0100010001010000_1;
      patterns[2120] = 17'b0000010010100001_0;
      patterns[2121] = 17'b1000010001010111_0;
      patterns[2122] = 17'b1001010001010111_0;
      patterns[2123] = 17'b1010010001010111_0;
      patterns[2124] = 17'b1011010001010111_0;
      patterns[2125] = 17'b0101010001010000_0;
      patterns[2126] = 17'b0100010001010000_1;
      patterns[2127] = 17'b0000010010101001_0;
      patterns[2128] = 17'b1000010001100000_0;
      patterns[2129] = 17'b1001010001100000_0;
      patterns[2130] = 17'b1010010001100000_0;
      patterns[2131] = 17'b1011010001100000_0;
      patterns[2132] = 17'b0101010001100000_0;
      patterns[2133] = 17'b0100010001100000_1;
      patterns[2134] = 17'b0000010010101001_0;
      patterns[2135] = 17'b1000010001100001_0;
      patterns[2136] = 17'b1001010001100001_0;
      patterns[2137] = 17'b1010010001100001_0;
      patterns[2138] = 17'b1011010001100001_0;
      patterns[2139] = 17'b0101010001100000_0;
      patterns[2140] = 17'b0100010001100000_1;
      patterns[2141] = 17'b0000010010110000_0;
      patterns[2142] = 17'b1000010001100010_0;
      patterns[2143] = 17'b1001010001100010_0;
      patterns[2144] = 17'b1010010001100010_0;
      patterns[2145] = 17'b1011010001100010_0;
      patterns[2146] = 17'b0101010001100000_0;
      patterns[2147] = 17'b0100010001100000_1;
      patterns[2148] = 17'b0000010001101010_0;
      patterns[2149] = 17'b1000010001100011_0;
      patterns[2150] = 17'b1001010001100011_0;
      patterns[2151] = 17'b1010010001100011_0;
      patterns[2152] = 17'b1011010001100011_0;
      patterns[2153] = 17'b0101010001100000_0;
      patterns[2154] = 17'b0100010001100000_1;
      patterns[2155] = 17'b0000010011001001_0;
      patterns[2156] = 17'b1000010001100100_0;
      patterns[2157] = 17'b1001010001100100_0;
      patterns[2158] = 17'b1010010001100100_0;
      patterns[2159] = 17'b1011010001100100_0;
      patterns[2160] = 17'b0101010001100000_0;
      patterns[2161] = 17'b0100010001100000_1;
      patterns[2162] = 17'b0000010011111010_0;
      patterns[2163] = 17'b1000010001100101_0;
      patterns[2164] = 17'b1001010001100101_0;
      patterns[2165] = 17'b1010010001100101_0;
      patterns[2166] = 17'b1011010001100101_0;
      patterns[2167] = 17'b0101010001100000_0;
      patterns[2168] = 17'b0100010001100000_1;
      patterns[2169] = 17'b0000010010100000_0;
      patterns[2170] = 17'b1000010001100110_0;
      patterns[2171] = 17'b1001010001100110_0;
      patterns[2172] = 17'b1010010001100110_0;
      patterns[2173] = 17'b1011010001100110_0;
      patterns[2174] = 17'b0101010001100000_0;
      patterns[2175] = 17'b0100010001100000_1;
      patterns[2176] = 17'b0000010000001011_0;
      patterns[2177] = 17'b1000010001100111_0;
      patterns[2178] = 17'b1001010001100111_0;
      patterns[2179] = 17'b1010010001100111_0;
      patterns[2180] = 17'b1011010001100111_0;
      patterns[2181] = 17'b0101010001100000_0;
      patterns[2182] = 17'b0100010001100000_1;
      patterns[2183] = 17'b0000010010100001_0;
      patterns[2184] = 17'b1000010001110000_0;
      patterns[2185] = 17'b1001010001110000_0;
      patterns[2186] = 17'b1010010001110000_0;
      patterns[2187] = 17'b1011010001110000_0;
      patterns[2188] = 17'b0101010001110000_0;
      patterns[2189] = 17'b0100010001110000_1;
      patterns[2190] = 17'b0000010001010001_0;
      patterns[2191] = 17'b1000010001110001_0;
      patterns[2192] = 17'b1001010001110001_0;
      patterns[2193] = 17'b1010010001110001_0;
      patterns[2194] = 17'b1011010001110001_0;
      patterns[2195] = 17'b0101010001110000_0;
      patterns[2196] = 17'b0100010001110000_1;
      patterns[2197] = 17'b0000010000110101_0;
      patterns[2198] = 17'b1000010001110010_0;
      patterns[2199] = 17'b1001010001110010_0;
      patterns[2200] = 17'b1010010001110010_0;
      patterns[2201] = 17'b1011010001110010_0;
      patterns[2202] = 17'b0101010001110000_0;
      patterns[2203] = 17'b0100010001110000_1;
      patterns[2204] = 17'b0000010001101111_0;
      patterns[2205] = 17'b1000010001110011_0;
      patterns[2206] = 17'b1001010001110011_0;
      patterns[2207] = 17'b1010010001110011_0;
      patterns[2208] = 17'b1011010001110011_0;
      patterns[2209] = 17'b0101010001110000_0;
      patterns[2210] = 17'b0100010001110000_1;
      patterns[2211] = 17'b0000010011101101_0;
      patterns[2212] = 17'b1000010001110100_0;
      patterns[2213] = 17'b1001010001110100_0;
      patterns[2214] = 17'b1010010001110100_0;
      patterns[2215] = 17'b1011010001110100_0;
      patterns[2216] = 17'b0101010001110000_0;
      patterns[2217] = 17'b0100010001110000_1;
      patterns[2218] = 17'b0000010000110010_0;
      patterns[2219] = 17'b1000010001110101_0;
      patterns[2220] = 17'b1001010001110101_0;
      patterns[2221] = 17'b1010010001110101_0;
      patterns[2222] = 17'b1011010001110101_0;
      patterns[2223] = 17'b0101010001110000_0;
      patterns[2224] = 17'b0100010001110000_1;
      patterns[2225] = 17'b0000010000110110_0;
      patterns[2226] = 17'b1000010001110110_0;
      patterns[2227] = 17'b1001010001110110_0;
      patterns[2228] = 17'b1010010001110110_0;
      patterns[2229] = 17'b1011010001110110_0;
      patterns[2230] = 17'b0101010001110000_0;
      patterns[2231] = 17'b0100010001110000_1;
      patterns[2232] = 17'b0000010011100010_0;
      patterns[2233] = 17'b1000010001110111_0;
      patterns[2234] = 17'b1001010001110111_0;
      patterns[2235] = 17'b1010010001110111_0;
      patterns[2236] = 17'b1011010001110111_0;
      patterns[2237] = 17'b0101010001110000_0;
      patterns[2238] = 17'b0100010001110000_1;
      patterns[2239] = 17'b0000010001000001_0;
      patterns[2240] = 17'b1000010100000000_0;
      patterns[2241] = 17'b1001010100000000_0;
      patterns[2242] = 17'b1010010100000000_0;
      patterns[2243] = 17'b1011010100000000_0;
      patterns[2244] = 17'b0101010100000000_0;
      patterns[2245] = 17'b0100010100000000_1;
      patterns[2246] = 17'b0000010111110011_0;
      patterns[2247] = 17'b1000010100000001_0;
      patterns[2248] = 17'b1001010100000001_0;
      patterns[2249] = 17'b1010010100000001_0;
      patterns[2250] = 17'b1011010100000001_0;
      patterns[2251] = 17'b0101010100000000_0;
      patterns[2252] = 17'b0100010100000000_1;
      patterns[2253] = 17'b0000010100011000_0;
      patterns[2254] = 17'b1000010100000010_0;
      patterns[2255] = 17'b1001010100000010_0;
      patterns[2256] = 17'b1010010100000010_0;
      patterns[2257] = 17'b1011010100000010_0;
      patterns[2258] = 17'b0101010100000000_0;
      patterns[2259] = 17'b0100010100000000_1;
      patterns[2260] = 17'b0000010101100101_0;
      patterns[2261] = 17'b1000010100000011_0;
      patterns[2262] = 17'b1001010100000011_0;
      patterns[2263] = 17'b1010010100000011_0;
      patterns[2264] = 17'b1011010100000011_0;
      patterns[2265] = 17'b0101010100000000_0;
      patterns[2266] = 17'b0100010100000000_1;
      patterns[2267] = 17'b0000010101100011_0;
      patterns[2268] = 17'b1000010100000100_0;
      patterns[2269] = 17'b1001010100000100_0;
      patterns[2270] = 17'b1010010100000100_0;
      patterns[2271] = 17'b1011010100000100_0;
      patterns[2272] = 17'b0101010100000000_0;
      patterns[2273] = 17'b0100010100000000_1;
      patterns[2274] = 17'b0000010100000101_0;
      patterns[2275] = 17'b1000010100000101_0;
      patterns[2276] = 17'b1001010100000101_0;
      patterns[2277] = 17'b1010010100000101_0;
      patterns[2278] = 17'b1011010100000101_0;
      patterns[2279] = 17'b0101010100000000_0;
      patterns[2280] = 17'b0100010100000000_1;
      patterns[2281] = 17'b0000010100111101_0;
      patterns[2282] = 17'b1000010100000110_0;
      patterns[2283] = 17'b1001010100000110_0;
      patterns[2284] = 17'b1010010100000110_0;
      patterns[2285] = 17'b1011010100000110_0;
      patterns[2286] = 17'b0101010100000000_0;
      patterns[2287] = 17'b0100010100000000_1;
      patterns[2288] = 17'b0000010110101000_0;
      patterns[2289] = 17'b1000010100000111_0;
      patterns[2290] = 17'b1001010100000111_0;
      patterns[2291] = 17'b1010010100000111_0;
      patterns[2292] = 17'b1011010100000111_0;
      patterns[2293] = 17'b0101010100000000_0;
      patterns[2294] = 17'b0100010100000000_1;
      patterns[2295] = 17'b0000010110101111_0;
      patterns[2296] = 17'b1000010100010000_0;
      patterns[2297] = 17'b1001010100010000_0;
      patterns[2298] = 17'b1010010100010000_0;
      patterns[2299] = 17'b1011010100010000_0;
      patterns[2300] = 17'b0101010100010000_0;
      patterns[2301] = 17'b0100010100010000_1;
      patterns[2302] = 17'b0000010111010010_0;
      patterns[2303] = 17'b1000010100010001_0;
      patterns[2304] = 17'b1001010100010001_0;
      patterns[2305] = 17'b1010010100010001_0;
      patterns[2306] = 17'b1011010100010001_0;
      patterns[2307] = 17'b0101010100010000_0;
      patterns[2308] = 17'b0100010100010000_1;
      patterns[2309] = 17'b0000010111010001_0;
      patterns[2310] = 17'b1000010100010010_0;
      patterns[2311] = 17'b1001010100010010_0;
      patterns[2312] = 17'b1010010100010010_0;
      patterns[2313] = 17'b1011010100010010_0;
      patterns[2314] = 17'b0101010100010000_0;
      patterns[2315] = 17'b0100010100010000_1;
      patterns[2316] = 17'b0000010101001010_0;
      patterns[2317] = 17'b1000010100010011_0;
      patterns[2318] = 17'b1001010100010011_0;
      patterns[2319] = 17'b1010010100010011_0;
      patterns[2320] = 17'b1011010100010011_0;
      patterns[2321] = 17'b0101010100010000_0;
      patterns[2322] = 17'b0100010100010000_1;
      patterns[2323] = 17'b0000010100010011_0;
      patterns[2324] = 17'b1000010100010100_0;
      patterns[2325] = 17'b1001010100010100_0;
      patterns[2326] = 17'b1010010100010100_0;
      patterns[2327] = 17'b1011010100010100_0;
      patterns[2328] = 17'b0101010100010000_0;
      patterns[2329] = 17'b0100010100010000_1;
      patterns[2330] = 17'b0000010111111010_0;
      patterns[2331] = 17'b1000010100010101_0;
      patterns[2332] = 17'b1001010100010101_0;
      patterns[2333] = 17'b1010010100010101_0;
      patterns[2334] = 17'b1011010100010101_0;
      patterns[2335] = 17'b0101010100010000_0;
      patterns[2336] = 17'b0100010100010000_1;
      patterns[2337] = 17'b0000010100011110_0;
      patterns[2338] = 17'b1000010100010110_0;
      patterns[2339] = 17'b1001010100010110_0;
      patterns[2340] = 17'b1010010100010110_0;
      patterns[2341] = 17'b1011010100010110_0;
      patterns[2342] = 17'b0101010100010000_0;
      patterns[2343] = 17'b0100010100010000_1;
      patterns[2344] = 17'b0000010111100111_0;
      patterns[2345] = 17'b1000010100010111_0;
      patterns[2346] = 17'b1001010100010111_0;
      patterns[2347] = 17'b1010010100010111_0;
      patterns[2348] = 17'b1011010100010111_0;
      patterns[2349] = 17'b0101010100010000_0;
      patterns[2350] = 17'b0100010100010000_1;
      patterns[2351] = 17'b0000010101100011_0;
      patterns[2352] = 17'b1000010100100000_0;
      patterns[2353] = 17'b1001010100100000_0;
      patterns[2354] = 17'b1010010100100000_0;
      patterns[2355] = 17'b1011010100100000_0;
      patterns[2356] = 17'b0101010100100000_0;
      patterns[2357] = 17'b0100010100100000_1;
      patterns[2358] = 17'b0000010111101001_0;
      patterns[2359] = 17'b1000010100100001_0;
      patterns[2360] = 17'b1001010100100001_0;
      patterns[2361] = 17'b1010010100100001_0;
      patterns[2362] = 17'b1011010100100001_0;
      patterns[2363] = 17'b0101010100100000_0;
      patterns[2364] = 17'b0100010100100000_1;
      patterns[2365] = 17'b0000010111101000_0;
      patterns[2366] = 17'b1000010100100010_0;
      patterns[2367] = 17'b1001010100100010_0;
      patterns[2368] = 17'b1010010100100010_0;
      patterns[2369] = 17'b1011010100100010_0;
      patterns[2370] = 17'b0101010100100000_0;
      patterns[2371] = 17'b0100010100100000_1;
      patterns[2372] = 17'b0000010111100001_0;
      patterns[2373] = 17'b1000010100100011_0;
      patterns[2374] = 17'b1001010100100011_0;
      patterns[2375] = 17'b1010010100100011_0;
      patterns[2376] = 17'b1011010100100011_0;
      patterns[2377] = 17'b0101010100100000_0;
      patterns[2378] = 17'b0100010100100000_1;
      patterns[2379] = 17'b0000010110010001_0;
      patterns[2380] = 17'b1000010100100100_0;
      patterns[2381] = 17'b1001010100100100_0;
      patterns[2382] = 17'b1010010100100100_0;
      patterns[2383] = 17'b1011010100100100_0;
      patterns[2384] = 17'b0101010100100000_0;
      patterns[2385] = 17'b0100010100100000_1;
      patterns[2386] = 17'b0000010101101010_0;
      patterns[2387] = 17'b1000010100100101_0;
      patterns[2388] = 17'b1001010100100101_0;
      patterns[2389] = 17'b1010010100100101_0;
      patterns[2390] = 17'b1011010100100101_0;
      patterns[2391] = 17'b0101010100100000_0;
      patterns[2392] = 17'b0100010100100000_1;
      patterns[2393] = 17'b0000010101111101_0;
      patterns[2394] = 17'b1000010100100110_0;
      patterns[2395] = 17'b1001010100100110_0;
      patterns[2396] = 17'b1010010100100110_0;
      patterns[2397] = 17'b1011010100100110_0;
      patterns[2398] = 17'b0101010100100000_0;
      patterns[2399] = 17'b0100010100100000_1;
      patterns[2400] = 17'b0000010101011101_0;
      patterns[2401] = 17'b1000010100100111_0;
      patterns[2402] = 17'b1001010100100111_0;
      patterns[2403] = 17'b1010010100100111_0;
      patterns[2404] = 17'b1011010100100111_0;
      patterns[2405] = 17'b0101010100100000_0;
      patterns[2406] = 17'b0100010100100000_1;
      patterns[2407] = 17'b0000010110101011_0;
      patterns[2408] = 17'b1000010100110000_0;
      patterns[2409] = 17'b1001010100110000_0;
      patterns[2410] = 17'b1010010100110000_0;
      patterns[2411] = 17'b1011010100110000_0;
      patterns[2412] = 17'b0101010100110000_0;
      patterns[2413] = 17'b0100010100110000_1;
      patterns[2414] = 17'b0000010110010110_0;
      patterns[2415] = 17'b1000010100110001_0;
      patterns[2416] = 17'b1001010100110001_0;
      patterns[2417] = 17'b1010010100110001_0;
      patterns[2418] = 17'b1011010100110001_0;
      patterns[2419] = 17'b0101010100110000_0;
      patterns[2420] = 17'b0100010100110000_1;
      patterns[2421] = 17'b0000010111100110_0;
      patterns[2422] = 17'b1000010100110010_0;
      patterns[2423] = 17'b1001010100110010_0;
      patterns[2424] = 17'b1010010100110010_0;
      patterns[2425] = 17'b1011010100110010_0;
      patterns[2426] = 17'b0101010100110000_0;
      patterns[2427] = 17'b0100010100110000_1;
      patterns[2428] = 17'b0000010111000110_0;
      patterns[2429] = 17'b1000010100110011_0;
      patterns[2430] = 17'b1001010100110011_0;
      patterns[2431] = 17'b1010010100110011_0;
      patterns[2432] = 17'b1011010100110011_0;
      patterns[2433] = 17'b0101010100110000_0;
      patterns[2434] = 17'b0100010100110000_1;
      patterns[2435] = 17'b0000010101001000_0;
      patterns[2436] = 17'b1000010100110100_0;
      patterns[2437] = 17'b1001010100110100_0;
      patterns[2438] = 17'b1010010100110100_0;
      patterns[2439] = 17'b1011010100110100_0;
      patterns[2440] = 17'b0101010100110000_0;
      patterns[2441] = 17'b0100010100110000_1;
      patterns[2442] = 17'b0000010110110101_0;
      patterns[2443] = 17'b1000010100110101_0;
      patterns[2444] = 17'b1001010100110101_0;
      patterns[2445] = 17'b1010010100110101_0;
      patterns[2446] = 17'b1011010100110101_0;
      patterns[2447] = 17'b0101010100110000_0;
      patterns[2448] = 17'b0100010100110000_1;
      patterns[2449] = 17'b0000010111001110_0;
      patterns[2450] = 17'b1000010100110110_0;
      patterns[2451] = 17'b1001010100110110_0;
      patterns[2452] = 17'b1010010100110110_0;
      patterns[2453] = 17'b1011010100110110_0;
      patterns[2454] = 17'b0101010100110000_0;
      patterns[2455] = 17'b0100010100110000_1;
      patterns[2456] = 17'b0000010101010000_0;
      patterns[2457] = 17'b1000010100110111_0;
      patterns[2458] = 17'b1001010100110111_0;
      patterns[2459] = 17'b1010010100110111_0;
      patterns[2460] = 17'b1011010100110111_0;
      patterns[2461] = 17'b0101010100110000_0;
      patterns[2462] = 17'b0100010100110000_1;
      patterns[2463] = 17'b0000010101110101_0;
      patterns[2464] = 17'b1000010101000000_0;
      patterns[2465] = 17'b1001010101000000_0;
      patterns[2466] = 17'b1010010101000000_0;
      patterns[2467] = 17'b1011010101000000_0;
      patterns[2468] = 17'b0101010101000000_0;
      patterns[2469] = 17'b0100010101000000_1;
      patterns[2470] = 17'b0000010100000111_0;
      patterns[2471] = 17'b1000010101000001_0;
      patterns[2472] = 17'b1001010101000001_0;
      patterns[2473] = 17'b1010010101000001_0;
      patterns[2474] = 17'b1011010101000001_0;
      patterns[2475] = 17'b0101010101000000_0;
      patterns[2476] = 17'b0100010101000000_1;
      patterns[2477] = 17'b0000010110001101_0;
      patterns[2478] = 17'b1000010101000010_0;
      patterns[2479] = 17'b1001010101000010_0;
      patterns[2480] = 17'b1010010101000010_0;
      patterns[2481] = 17'b1011010101000010_0;
      patterns[2482] = 17'b0101010101000000_0;
      patterns[2483] = 17'b0100010101000000_1;
      patterns[2484] = 17'b0000010101011101_0;
      patterns[2485] = 17'b1000010101000011_0;
      patterns[2486] = 17'b1001010101000011_0;
      patterns[2487] = 17'b1010010101000011_0;
      patterns[2488] = 17'b1011010101000011_0;
      patterns[2489] = 17'b0101010101000000_0;
      patterns[2490] = 17'b0100010101000000_1;
      patterns[2491] = 17'b0000010100011010_0;
      patterns[2492] = 17'b1000010101000100_0;
      patterns[2493] = 17'b1001010101000100_0;
      patterns[2494] = 17'b1010010101000100_0;
      patterns[2495] = 17'b1011010101000100_0;
      patterns[2496] = 17'b0101010101000000_0;
      patterns[2497] = 17'b0100010101000000_1;
      patterns[2498] = 17'b0000010100011000_0;
      patterns[2499] = 17'b1000010101000101_0;
      patterns[2500] = 17'b1001010101000101_0;
      patterns[2501] = 17'b1010010101000101_0;
      patterns[2502] = 17'b1011010101000101_0;
      patterns[2503] = 17'b0101010101000000_0;
      patterns[2504] = 17'b0100010101000000_1;
      patterns[2505] = 17'b0000010111110011_0;
      patterns[2506] = 17'b1000010101000110_0;
      patterns[2507] = 17'b1001010101000110_0;
      patterns[2508] = 17'b1010010101000110_0;
      patterns[2509] = 17'b1011010101000110_0;
      patterns[2510] = 17'b0101010101000000_0;
      patterns[2511] = 17'b0100010101000000_1;
      patterns[2512] = 17'b0000010101100100_0;
      patterns[2513] = 17'b1000010101000111_0;
      patterns[2514] = 17'b1001010101000111_0;
      patterns[2515] = 17'b1010010101000111_0;
      patterns[2516] = 17'b1011010101000111_0;
      patterns[2517] = 17'b0101010101000000_0;
      patterns[2518] = 17'b0100010101000000_1;
      patterns[2519] = 17'b0000010100111111_0;
      patterns[2520] = 17'b1000010101010000_0;
      patterns[2521] = 17'b1001010101010000_0;
      patterns[2522] = 17'b1010010101010000_0;
      patterns[2523] = 17'b1011010101010000_0;
      patterns[2524] = 17'b0101010101010000_0;
      patterns[2525] = 17'b0100010101010000_1;
      patterns[2526] = 17'b0000010100111100_0;
      patterns[2527] = 17'b1000010101010001_0;
      patterns[2528] = 17'b1001010101010001_0;
      patterns[2529] = 17'b1010010101010001_0;
      patterns[2530] = 17'b1011010101010001_0;
      patterns[2531] = 17'b0101010101010000_0;
      patterns[2532] = 17'b0100010101010000_1;
      patterns[2533] = 17'b0000010101100001_0;
      patterns[2534] = 17'b1000010101010010_0;
      patterns[2535] = 17'b1001010101010010_0;
      patterns[2536] = 17'b1010010101010010_0;
      patterns[2537] = 17'b1011010101010010_0;
      patterns[2538] = 17'b0101010101010000_0;
      patterns[2539] = 17'b0100010101010000_1;
      patterns[2540] = 17'b0000010111101100_0;
      patterns[2541] = 17'b1000010101010011_0;
      patterns[2542] = 17'b1001010101010011_0;
      patterns[2543] = 17'b1010010101010011_0;
      patterns[2544] = 17'b1011010101010011_0;
      patterns[2545] = 17'b0101010101010000_0;
      patterns[2546] = 17'b0100010101010000_1;
      patterns[2547] = 17'b0000010101111100_0;
      patterns[2548] = 17'b1000010101010100_0;
      patterns[2549] = 17'b1001010101010100_0;
      patterns[2550] = 17'b1010010101010100_0;
      patterns[2551] = 17'b1011010101010100_0;
      patterns[2552] = 17'b0101010101010000_0;
      patterns[2553] = 17'b0100010101010000_1;
      patterns[2554] = 17'b0000010100100001_0;
      patterns[2555] = 17'b1000010101010101_0;
      patterns[2556] = 17'b1001010101010101_0;
      patterns[2557] = 17'b1010010101010101_0;
      patterns[2558] = 17'b1011010101010101_0;
      patterns[2559] = 17'b0101010101010000_0;
      patterns[2560] = 17'b0100010101010000_1;
      patterns[2561] = 17'b0000010111111010_0;
      patterns[2562] = 17'b1000010101010110_0;
      patterns[2563] = 17'b1001010101010110_0;
      patterns[2564] = 17'b1010010101010110_0;
      patterns[2565] = 17'b1011010101010110_0;
      patterns[2566] = 17'b0101010101010000_0;
      patterns[2567] = 17'b0100010101010000_1;
      patterns[2568] = 17'b0000010101110000_0;
      patterns[2569] = 17'b1000010101010111_0;
      patterns[2570] = 17'b1001010101010111_0;
      patterns[2571] = 17'b1010010101010111_0;
      patterns[2572] = 17'b1011010101010111_0;
      patterns[2573] = 17'b0101010101010000_0;
      patterns[2574] = 17'b0100010101010000_1;
      patterns[2575] = 17'b0000010101111100_0;
      patterns[2576] = 17'b1000010101100000_0;
      patterns[2577] = 17'b1001010101100000_0;
      patterns[2578] = 17'b1010010101100000_0;
      patterns[2579] = 17'b1011010101100000_0;
      patterns[2580] = 17'b0101010101100000_0;
      patterns[2581] = 17'b0100010101100000_1;
      patterns[2582] = 17'b0000010110111011_0;
      patterns[2583] = 17'b1000010101100001_0;
      patterns[2584] = 17'b1001010101100001_0;
      patterns[2585] = 17'b1010010101100001_0;
      patterns[2586] = 17'b1011010101100001_0;
      patterns[2587] = 17'b0101010101100000_0;
      patterns[2588] = 17'b0100010101100000_1;
      patterns[2589] = 17'b0000010110110100_0;
      patterns[2590] = 17'b1000010101100010_0;
      patterns[2591] = 17'b1001010101100010_0;
      patterns[2592] = 17'b1010010101100010_0;
      patterns[2593] = 17'b1011010101100010_0;
      patterns[2594] = 17'b0101010101100000_0;
      patterns[2595] = 17'b0100010101100000_1;
      patterns[2596] = 17'b0000010110011101_0;
      patterns[2597] = 17'b1000010101100011_0;
      patterns[2598] = 17'b1001010101100011_0;
      patterns[2599] = 17'b1010010101100011_0;
      patterns[2600] = 17'b1011010101100011_0;
      patterns[2601] = 17'b0101010101100000_0;
      patterns[2602] = 17'b0100010101100000_1;
      patterns[2603] = 17'b0000010101101100_0;
      patterns[2604] = 17'b1000010101100100_0;
      patterns[2605] = 17'b1001010101100100_0;
      patterns[2606] = 17'b1010010101100100_0;
      patterns[2607] = 17'b1011010101100100_0;
      patterns[2608] = 17'b0101010101100000_0;
      patterns[2609] = 17'b0100010101100000_1;
      patterns[2610] = 17'b0000010111110110_0;
      patterns[2611] = 17'b1000010101100101_0;
      patterns[2612] = 17'b1001010101100101_0;
      patterns[2613] = 17'b1010010101100101_0;
      patterns[2614] = 17'b1011010101100101_0;
      patterns[2615] = 17'b0101010101100000_0;
      patterns[2616] = 17'b0100010101100000_1;
      patterns[2617] = 17'b0000010101011101_0;
      patterns[2618] = 17'b1000010101100110_0;
      patterns[2619] = 17'b1001010101100110_0;
      patterns[2620] = 17'b1010010101100110_0;
      patterns[2621] = 17'b1011010101100110_0;
      patterns[2622] = 17'b0101010101100000_0;
      patterns[2623] = 17'b0100010101100000_1;
      patterns[2624] = 17'b0000010100011101_0;
      patterns[2625] = 17'b1000010101100111_0;
      patterns[2626] = 17'b1001010101100111_0;
      patterns[2627] = 17'b1010010101100111_0;
      patterns[2628] = 17'b1011010101100111_0;
      patterns[2629] = 17'b0101010101100000_0;
      patterns[2630] = 17'b0100010101100000_1;
      patterns[2631] = 17'b0000010111000001_0;
      patterns[2632] = 17'b1000010101110000_0;
      patterns[2633] = 17'b1001010101110000_0;
      patterns[2634] = 17'b1010010101110000_0;
      patterns[2635] = 17'b1011010101110000_0;
      patterns[2636] = 17'b0101010101110000_0;
      patterns[2637] = 17'b0100010101110000_1;
      patterns[2638] = 17'b0000010101000011_0;
      patterns[2639] = 17'b1000010101110001_0;
      patterns[2640] = 17'b1001010101110001_0;
      patterns[2641] = 17'b1010010101110001_0;
      patterns[2642] = 17'b1011010101110001_0;
      patterns[2643] = 17'b0101010101110000_0;
      patterns[2644] = 17'b0100010101110000_1;
      patterns[2645] = 17'b0000010111000011_0;
      patterns[2646] = 17'b1000010101110010_0;
      patterns[2647] = 17'b1001010101110010_0;
      patterns[2648] = 17'b1010010101110010_0;
      patterns[2649] = 17'b1011010101110010_0;
      patterns[2650] = 17'b0101010101110000_0;
      patterns[2651] = 17'b0100010101110000_1;
      patterns[2652] = 17'b0000010101000100_0;
      patterns[2653] = 17'b1000010101110011_0;
      patterns[2654] = 17'b1001010101110011_0;
      patterns[2655] = 17'b1010010101110011_0;
      patterns[2656] = 17'b1011010101110011_0;
      patterns[2657] = 17'b0101010101110000_0;
      patterns[2658] = 17'b0100010101110000_1;
      patterns[2659] = 17'b0000010111010011_0;
      patterns[2660] = 17'b1000010101110100_0;
      patterns[2661] = 17'b1001010101110100_0;
      patterns[2662] = 17'b1010010101110100_0;
      patterns[2663] = 17'b1011010101110100_0;
      patterns[2664] = 17'b0101010101110000_0;
      patterns[2665] = 17'b0100010101110000_1;
      patterns[2666] = 17'b0000010111100110_0;
      patterns[2667] = 17'b1000010101110101_0;
      patterns[2668] = 17'b1001010101110101_0;
      patterns[2669] = 17'b1010010101110101_0;
      patterns[2670] = 17'b1011010101110101_0;
      patterns[2671] = 17'b0101010101110000_0;
      patterns[2672] = 17'b0100010101110000_1;
      patterns[2673] = 17'b0000010101101011_0;
      patterns[2674] = 17'b1000010101110110_0;
      patterns[2675] = 17'b1001010101110110_0;
      patterns[2676] = 17'b1010010101110110_0;
      patterns[2677] = 17'b1011010101110110_0;
      patterns[2678] = 17'b0101010101110000_0;
      patterns[2679] = 17'b0100010101110000_1;
      patterns[2680] = 17'b0000010101100001_0;
      patterns[2681] = 17'b1000010101110111_0;
      patterns[2682] = 17'b1001010101110111_0;
      patterns[2683] = 17'b1010010101110111_0;
      patterns[2684] = 17'b1011010101110111_0;
      patterns[2685] = 17'b0101010101110000_0;
      patterns[2686] = 17'b0100010101110000_1;
      patterns[2687] = 17'b0000010110000010_0;
      patterns[2688] = 17'b1000011000000000_0;
      patterns[2689] = 17'b1001011000000000_0;
      patterns[2690] = 17'b1010011000000000_0;
      patterns[2691] = 17'b1011011000000000_0;
      patterns[2692] = 17'b0101011000000000_0;
      patterns[2693] = 17'b0100011000000000_1;
      patterns[2694] = 17'b0000011000101101_0;
      patterns[2695] = 17'b1000011000000001_0;
      patterns[2696] = 17'b1001011000000001_0;
      patterns[2697] = 17'b1010011000000001_0;
      patterns[2698] = 17'b1011011000000001_0;
      patterns[2699] = 17'b0101011000000000_0;
      patterns[2700] = 17'b0100011000000000_1;
      patterns[2701] = 17'b0000011010011110_0;
      patterns[2702] = 17'b1000011000000010_0;
      patterns[2703] = 17'b1001011000000010_0;
      patterns[2704] = 17'b1010011000000010_0;
      patterns[2705] = 17'b1011011000000010_0;
      patterns[2706] = 17'b0101011000000000_0;
      patterns[2707] = 17'b0100011000000000_1;
      patterns[2708] = 17'b0000011000010110_0;
      patterns[2709] = 17'b1000011000000011_0;
      patterns[2710] = 17'b1001011000000011_0;
      patterns[2711] = 17'b1010011000000011_0;
      patterns[2712] = 17'b1011011000000011_0;
      patterns[2713] = 17'b0101011000000000_0;
      patterns[2714] = 17'b0100011000000000_1;
      patterns[2715] = 17'b0000011000010001_0;
      patterns[2716] = 17'b1000011000000100_0;
      patterns[2717] = 17'b1001011000000100_0;
      patterns[2718] = 17'b1010011000000100_0;
      patterns[2719] = 17'b1011011000000100_0;
      patterns[2720] = 17'b0101011000000000_0;
      patterns[2721] = 17'b0100011000000000_1;
      patterns[2722] = 17'b0000011000000100_0;
      patterns[2723] = 17'b1000011000000101_0;
      patterns[2724] = 17'b1001011000000101_0;
      patterns[2725] = 17'b1010011000000101_0;
      patterns[2726] = 17'b1011011000000101_0;
      patterns[2727] = 17'b0101011000000000_0;
      patterns[2728] = 17'b0100011000000000_1;
      patterns[2729] = 17'b0000011010101110_0;
      patterns[2730] = 17'b1000011000000110_0;
      patterns[2731] = 17'b1001011000000110_0;
      patterns[2732] = 17'b1010011000000110_0;
      patterns[2733] = 17'b1011011000000110_0;
      patterns[2734] = 17'b0101011000000000_0;
      patterns[2735] = 17'b0100011000000000_1;
      patterns[2736] = 17'b0000011000010000_0;
      patterns[2737] = 17'b1000011000000111_0;
      patterns[2738] = 17'b1001011000000111_0;
      patterns[2739] = 17'b1010011000000111_0;
      patterns[2740] = 17'b1011011000000111_0;
      patterns[2741] = 17'b0101011000000000_0;
      patterns[2742] = 17'b0100011000000000_1;
      patterns[2743] = 17'b0000011001000011_0;
      patterns[2744] = 17'b1000011000010000_0;
      patterns[2745] = 17'b1001011000010000_0;
      patterns[2746] = 17'b1010011000010000_0;
      patterns[2747] = 17'b1011011000010000_0;
      patterns[2748] = 17'b0101011000010000_0;
      patterns[2749] = 17'b0100011000010000_1;
      patterns[2750] = 17'b0000011000111111_0;
      patterns[2751] = 17'b1000011000010001_0;
      patterns[2752] = 17'b1001011000010001_0;
      patterns[2753] = 17'b1010011000010001_0;
      patterns[2754] = 17'b1011011000010001_0;
      patterns[2755] = 17'b0101011000010000_0;
      patterns[2756] = 17'b0100011000010000_1;
      patterns[2757] = 17'b0000011011011101_0;
      patterns[2758] = 17'b1000011000010010_0;
      patterns[2759] = 17'b1001011000010010_0;
      patterns[2760] = 17'b1010011000010010_0;
      patterns[2761] = 17'b1011011000010010_0;
      patterns[2762] = 17'b0101011000010000_0;
      patterns[2763] = 17'b0100011000010000_1;
      patterns[2764] = 17'b0000011010111101_0;
      patterns[2765] = 17'b1000011000010011_0;
      patterns[2766] = 17'b1001011000010011_0;
      patterns[2767] = 17'b1010011000010011_0;
      patterns[2768] = 17'b1011011000010011_0;
      patterns[2769] = 17'b0101011000010000_0;
      patterns[2770] = 17'b0100011000010000_1;
      patterns[2771] = 17'b0000011011011011_0;
      patterns[2772] = 17'b1000011000010100_0;
      patterns[2773] = 17'b1001011000010100_0;
      patterns[2774] = 17'b1010011000010100_0;
      patterns[2775] = 17'b1011011000010100_0;
      patterns[2776] = 17'b0101011000010000_0;
      patterns[2777] = 17'b0100011000010000_1;
      patterns[2778] = 17'b0000011010111101_0;
      patterns[2779] = 17'b1000011000010101_0;
      patterns[2780] = 17'b1001011000010101_0;
      patterns[2781] = 17'b1010011000010101_0;
      patterns[2782] = 17'b1011011000010101_0;
      patterns[2783] = 17'b0101011000010000_0;
      patterns[2784] = 17'b0100011000010000_1;
      patterns[2785] = 17'b0000011001111111_0;
      patterns[2786] = 17'b1000011000010110_0;
      patterns[2787] = 17'b1001011000010110_0;
      patterns[2788] = 17'b1010011000010110_0;
      patterns[2789] = 17'b1011011000010110_0;
      patterns[2790] = 17'b0101011000010000_0;
      patterns[2791] = 17'b0100011000010000_1;
      patterns[2792] = 17'b0000011000010111_0;
      patterns[2793] = 17'b1000011000010111_0;
      patterns[2794] = 17'b1001011000010111_0;
      patterns[2795] = 17'b1010011000010111_0;
      patterns[2796] = 17'b1011011000010111_0;
      patterns[2797] = 17'b0101011000010000_0;
      patterns[2798] = 17'b0100011000010000_1;
      patterns[2799] = 17'b0000011001101110_0;
      patterns[2800] = 17'b1000011000100000_0;
      patterns[2801] = 17'b1001011000100000_0;
      patterns[2802] = 17'b1010011000100000_0;
      patterns[2803] = 17'b1011011000100000_0;
      patterns[2804] = 17'b0101011000100000_0;
      patterns[2805] = 17'b0100011000100000_1;
      patterns[2806] = 17'b0000011000010010_0;
      patterns[2807] = 17'b1000011000100001_0;
      patterns[2808] = 17'b1001011000100001_0;
      patterns[2809] = 17'b1010011000100001_0;
      patterns[2810] = 17'b1011011000100001_0;
      patterns[2811] = 17'b0101011000100000_0;
      patterns[2812] = 17'b0100011000100000_1;
      patterns[2813] = 17'b0000011001101000_0;
      patterns[2814] = 17'b1000011000100010_0;
      patterns[2815] = 17'b1001011000100010_0;
      patterns[2816] = 17'b1010011000100010_0;
      patterns[2817] = 17'b1011011000100010_0;
      patterns[2818] = 17'b0101011000100000_0;
      patterns[2819] = 17'b0100011000100000_1;
      patterns[2820] = 17'b0000011001101111_0;
      patterns[2821] = 17'b1000011000100011_0;
      patterns[2822] = 17'b1001011000100011_0;
      patterns[2823] = 17'b1010011000100011_0;
      patterns[2824] = 17'b1011011000100011_0;
      patterns[2825] = 17'b0101011000100000_0;
      patterns[2826] = 17'b0100011000100000_1;
      patterns[2827] = 17'b0000011010110001_0;
      patterns[2828] = 17'b1000011000100100_0;
      patterns[2829] = 17'b1001011000100100_0;
      patterns[2830] = 17'b1010011000100100_0;
      patterns[2831] = 17'b1011011000100100_0;
      patterns[2832] = 17'b0101011000100000_0;
      patterns[2833] = 17'b0100011000100000_1;
      patterns[2834] = 17'b0000011010100111_0;
      patterns[2835] = 17'b1000011000100101_0;
      patterns[2836] = 17'b1001011000100101_0;
      patterns[2837] = 17'b1010011000100101_0;
      patterns[2838] = 17'b1011011000100101_0;
      patterns[2839] = 17'b0101011000100000_0;
      patterns[2840] = 17'b0100011000100000_1;
      patterns[2841] = 17'b0000011000100001_0;
      patterns[2842] = 17'b1000011000100110_0;
      patterns[2843] = 17'b1001011000100110_0;
      patterns[2844] = 17'b1010011000100110_0;
      patterns[2845] = 17'b1011011000100110_0;
      patterns[2846] = 17'b0101011000100000_0;
      patterns[2847] = 17'b0100011000100000_1;
      patterns[2848] = 17'b0000011000101101_0;
      patterns[2849] = 17'b1000011000100111_0;
      patterns[2850] = 17'b1001011000100111_0;
      patterns[2851] = 17'b1010011000100111_0;
      patterns[2852] = 17'b1011011000100111_0;
      patterns[2853] = 17'b0101011000100000_0;
      patterns[2854] = 17'b0100011000100000_1;
      patterns[2855] = 17'b0000011001001011_0;
      patterns[2856] = 17'b1000011000110000_0;
      patterns[2857] = 17'b1001011000110000_0;
      patterns[2858] = 17'b1010011000110000_0;
      patterns[2859] = 17'b1011011000110000_0;
      patterns[2860] = 17'b0101011000110000_0;
      patterns[2861] = 17'b0100011000110000_1;
      patterns[2862] = 17'b0000011001101010_0;
      patterns[2863] = 17'b1000011000110001_0;
      patterns[2864] = 17'b1001011000110001_0;
      patterns[2865] = 17'b1010011000110001_0;
      patterns[2866] = 17'b1011011000110001_0;
      patterns[2867] = 17'b0101011000110000_0;
      patterns[2868] = 17'b0100011000110000_1;
      patterns[2869] = 17'b0000011011000111_0;
      patterns[2870] = 17'b1000011000110010_0;
      patterns[2871] = 17'b1001011000110010_0;
      patterns[2872] = 17'b1010011000110010_0;
      patterns[2873] = 17'b1011011000110010_0;
      patterns[2874] = 17'b0101011000110000_0;
      patterns[2875] = 17'b0100011000110000_1;
      patterns[2876] = 17'b0000011011110000_0;
      patterns[2877] = 17'b1000011000110011_0;
      patterns[2878] = 17'b1001011000110011_0;
      patterns[2879] = 17'b1010011000110011_0;
      patterns[2880] = 17'b1011011000110011_0;
      patterns[2881] = 17'b0101011000110000_0;
      patterns[2882] = 17'b0100011000110000_1;
      patterns[2883] = 17'b0000011001111001_0;
      patterns[2884] = 17'b1000011000110100_0;
      patterns[2885] = 17'b1001011000110100_0;
      patterns[2886] = 17'b1010011000110100_0;
      patterns[2887] = 17'b1011011000110100_0;
      patterns[2888] = 17'b0101011000110000_0;
      patterns[2889] = 17'b0100011000110000_1;
      patterns[2890] = 17'b0000011000000001_0;
      patterns[2891] = 17'b1000011000110101_0;
      patterns[2892] = 17'b1001011000110101_0;
      patterns[2893] = 17'b1010011000110101_0;
      patterns[2894] = 17'b1011011000110101_0;
      patterns[2895] = 17'b0101011000110000_0;
      patterns[2896] = 17'b0100011000110000_1;
      patterns[2897] = 17'b0000011011111101_0;
      patterns[2898] = 17'b1000011000110110_0;
      patterns[2899] = 17'b1001011000110110_0;
      patterns[2900] = 17'b1010011000110110_0;
      patterns[2901] = 17'b1011011000110110_0;
      patterns[2902] = 17'b0101011000110000_0;
      patterns[2903] = 17'b0100011000110000_1;
      patterns[2904] = 17'b0000011011110010_0;
      patterns[2905] = 17'b1000011000110111_0;
      patterns[2906] = 17'b1001011000110111_0;
      patterns[2907] = 17'b1010011000110111_0;
      patterns[2908] = 17'b1011011000110111_0;
      patterns[2909] = 17'b0101011000110000_0;
      patterns[2910] = 17'b0100011000110000_1;
      patterns[2911] = 17'b0000011010111011_0;
      patterns[2912] = 17'b1000011001000000_0;
      patterns[2913] = 17'b1001011001000000_0;
      patterns[2914] = 17'b1010011001000000_0;
      patterns[2915] = 17'b1011011001000000_0;
      patterns[2916] = 17'b0101011001000000_0;
      patterns[2917] = 17'b0100011001000000_1;
      patterns[2918] = 17'b0000011000001111_0;
      patterns[2919] = 17'b1000011001000001_0;
      patterns[2920] = 17'b1001011001000001_0;
      patterns[2921] = 17'b1010011001000001_0;
      patterns[2922] = 17'b1011011001000001_0;
      patterns[2923] = 17'b0101011001000000_0;
      patterns[2924] = 17'b0100011001000000_1;
      patterns[2925] = 17'b0000011011001110_0;
      patterns[2926] = 17'b1000011001000010_0;
      patterns[2927] = 17'b1001011001000010_0;
      patterns[2928] = 17'b1010011001000010_0;
      patterns[2929] = 17'b1011011001000010_0;
      patterns[2930] = 17'b0101011001000000_0;
      patterns[2931] = 17'b0100011001000000_1;
      patterns[2932] = 17'b0000011010101110_0;
      patterns[2933] = 17'b1000011001000011_0;
      patterns[2934] = 17'b1001011001000011_0;
      patterns[2935] = 17'b1010011001000011_0;
      patterns[2936] = 17'b1011011001000011_0;
      patterns[2937] = 17'b0101011001000000_0;
      patterns[2938] = 17'b0100011001000000_1;
      patterns[2939] = 17'b0000011000011101_0;
      patterns[2940] = 17'b1000011001000100_0;
      patterns[2941] = 17'b1001011001000100_0;
      patterns[2942] = 17'b1010011001000100_0;
      patterns[2943] = 17'b1011011001000100_0;
      patterns[2944] = 17'b0101011001000000_0;
      patterns[2945] = 17'b0100011001000000_1;
      patterns[2946] = 17'b0000011010100001_0;
      patterns[2947] = 17'b1000011001000101_0;
      patterns[2948] = 17'b1001011001000101_0;
      patterns[2949] = 17'b1010011001000101_0;
      patterns[2950] = 17'b1011011001000101_0;
      patterns[2951] = 17'b0101011001000000_0;
      patterns[2952] = 17'b0100011001000000_1;
      patterns[2953] = 17'b0000011011110100_0;
      patterns[2954] = 17'b1000011001000110_0;
      patterns[2955] = 17'b1001011001000110_0;
      patterns[2956] = 17'b1010011001000110_0;
      patterns[2957] = 17'b1011011001000110_0;
      patterns[2958] = 17'b0101011001000000_0;
      patterns[2959] = 17'b0100011001000000_1;
      patterns[2960] = 17'b0000011011011000_0;
      patterns[2961] = 17'b1000011001000111_0;
      patterns[2962] = 17'b1001011001000111_0;
      patterns[2963] = 17'b1010011001000111_0;
      patterns[2964] = 17'b1011011001000111_0;
      patterns[2965] = 17'b0101011001000000_0;
      patterns[2966] = 17'b0100011001000000_1;
      patterns[2967] = 17'b0000011010110011_0;
      patterns[2968] = 17'b1000011001010000_0;
      patterns[2969] = 17'b1001011001010000_0;
      patterns[2970] = 17'b1010011001010000_0;
      patterns[2971] = 17'b1011011001010000_0;
      patterns[2972] = 17'b0101011001010000_0;
      patterns[2973] = 17'b0100011001010000_1;
      patterns[2974] = 17'b0000011000000010_0;
      patterns[2975] = 17'b1000011001010001_0;
      patterns[2976] = 17'b1001011001010001_0;
      patterns[2977] = 17'b1010011001010001_0;
      patterns[2978] = 17'b1011011001010001_0;
      patterns[2979] = 17'b0101011001010000_0;
      patterns[2980] = 17'b0100011001010000_1;
      patterns[2981] = 17'b0000011010001101_0;
      patterns[2982] = 17'b1000011001010010_0;
      patterns[2983] = 17'b1001011001010010_0;
      patterns[2984] = 17'b1010011001010010_0;
      patterns[2985] = 17'b1011011001010010_0;
      patterns[2986] = 17'b0101011001010000_0;
      patterns[2987] = 17'b0100011001010000_1;
      patterns[2988] = 17'b0000011001010000_0;
      patterns[2989] = 17'b1000011001010011_0;
      patterns[2990] = 17'b1001011001010011_0;
      patterns[2991] = 17'b1010011001010011_0;
      patterns[2992] = 17'b1011011001010011_0;
      patterns[2993] = 17'b0101011001010000_0;
      patterns[2994] = 17'b0100011001010000_1;
      patterns[2995] = 17'b0000011000101110_0;
      patterns[2996] = 17'b1000011001010100_0;
      patterns[2997] = 17'b1001011001010100_0;
      patterns[2998] = 17'b1010011001010100_0;
      patterns[2999] = 17'b1011011001010100_0;
      patterns[3000] = 17'b0101011001010000_0;
      patterns[3001] = 17'b0100011001010000_1;
      patterns[3002] = 17'b0000011000111001_0;
      patterns[3003] = 17'b1000011001010101_0;
      patterns[3004] = 17'b1001011001010101_0;
      patterns[3005] = 17'b1010011001010101_0;
      patterns[3006] = 17'b1011011001010101_0;
      patterns[3007] = 17'b0101011001010000_0;
      patterns[3008] = 17'b0100011001010000_1;
      patterns[3009] = 17'b0000011011001011_0;
      patterns[3010] = 17'b1000011001010110_0;
      patterns[3011] = 17'b1001011001010110_0;
      patterns[3012] = 17'b1010011001010110_0;
      patterns[3013] = 17'b1011011001010110_0;
      patterns[3014] = 17'b0101011001010000_0;
      patterns[3015] = 17'b0100011001010000_1;
      patterns[3016] = 17'b0000011001010110_0;
      patterns[3017] = 17'b1000011001010111_0;
      patterns[3018] = 17'b1001011001010111_0;
      patterns[3019] = 17'b1010011001010111_0;
      patterns[3020] = 17'b1011011001010111_0;
      patterns[3021] = 17'b0101011001010000_0;
      patterns[3022] = 17'b0100011001010000_1;
      patterns[3023] = 17'b0000011010100001_0;
      patterns[3024] = 17'b1000011001100000_0;
      patterns[3025] = 17'b1001011001100000_0;
      patterns[3026] = 17'b1010011001100000_0;
      patterns[3027] = 17'b1011011001100000_0;
      patterns[3028] = 17'b0101011001100000_0;
      patterns[3029] = 17'b0100011001100000_1;
      patterns[3030] = 17'b0000011000110010_0;
      patterns[3031] = 17'b1000011001100001_0;
      patterns[3032] = 17'b1001011001100001_0;
      patterns[3033] = 17'b1010011001100001_0;
      patterns[3034] = 17'b1011011001100001_0;
      patterns[3035] = 17'b0101011001100000_0;
      patterns[3036] = 17'b0100011001100000_1;
      patterns[3037] = 17'b0000011011100100_0;
      patterns[3038] = 17'b1000011001100010_0;
      patterns[3039] = 17'b1001011001100010_0;
      patterns[3040] = 17'b1010011001100010_0;
      patterns[3041] = 17'b1011011001100010_0;
      patterns[3042] = 17'b0101011001100000_0;
      patterns[3043] = 17'b0100011001100000_1;
      patterns[3044] = 17'b0000011010000000_0;
      patterns[3045] = 17'b1000011001100011_0;
      patterns[3046] = 17'b1001011001100011_0;
      patterns[3047] = 17'b1010011001100011_0;
      patterns[3048] = 17'b1011011001100011_0;
      patterns[3049] = 17'b0101011001100000_0;
      patterns[3050] = 17'b0100011001100000_1;
      patterns[3051] = 17'b0000011011100110_0;
      patterns[3052] = 17'b1000011001100100_0;
      patterns[3053] = 17'b1001011001100100_0;
      patterns[3054] = 17'b1010011001100100_0;
      patterns[3055] = 17'b1011011001100100_0;
      patterns[3056] = 17'b0101011001100000_0;
      patterns[3057] = 17'b0100011001100000_1;
      patterns[3058] = 17'b0000011001000110_0;
      patterns[3059] = 17'b1000011001100101_0;
      patterns[3060] = 17'b1001011001100101_0;
      patterns[3061] = 17'b1010011001100101_0;
      patterns[3062] = 17'b1011011001100101_0;
      patterns[3063] = 17'b0101011001100000_0;
      patterns[3064] = 17'b0100011001100000_1;
      patterns[3065] = 17'b0000011000110100_0;
      patterns[3066] = 17'b1000011001100110_0;
      patterns[3067] = 17'b1001011001100110_0;
      patterns[3068] = 17'b1010011001100110_0;
      patterns[3069] = 17'b1011011001100110_0;
      patterns[3070] = 17'b0101011001100000_0;
      patterns[3071] = 17'b0100011001100000_1;
      patterns[3072] = 17'b0000011000101001_0;
      patterns[3073] = 17'b1000011001100111_0;
      patterns[3074] = 17'b1001011001100111_0;
      patterns[3075] = 17'b1010011001100111_0;
      patterns[3076] = 17'b1011011001100111_0;
      patterns[3077] = 17'b0101011001100000_0;
      patterns[3078] = 17'b0100011001100000_1;
      patterns[3079] = 17'b0000011000110011_0;
      patterns[3080] = 17'b1000011001110000_0;
      patterns[3081] = 17'b1001011001110000_0;
      patterns[3082] = 17'b1010011001110000_0;
      patterns[3083] = 17'b1011011001110000_0;
      patterns[3084] = 17'b0101011001110000_0;
      patterns[3085] = 17'b0100011001110000_1;
      patterns[3086] = 17'b0000011011110111_0;
      patterns[3087] = 17'b1000011001110001_0;
      patterns[3088] = 17'b1001011001110001_0;
      patterns[3089] = 17'b1010011001110001_0;
      patterns[3090] = 17'b1011011001110001_0;
      patterns[3091] = 17'b0101011001110000_0;
      patterns[3092] = 17'b0100011001110000_1;
      patterns[3093] = 17'b0000011000011001_0;
      patterns[3094] = 17'b1000011001110010_0;
      patterns[3095] = 17'b1001011001110010_0;
      patterns[3096] = 17'b1010011001110010_0;
      patterns[3097] = 17'b1011011001110010_0;
      patterns[3098] = 17'b0101011001110000_0;
      patterns[3099] = 17'b0100011001110000_1;
      patterns[3100] = 17'b0000011010101110_0;
      patterns[3101] = 17'b1000011001110011_0;
      patterns[3102] = 17'b1001011001110011_0;
      patterns[3103] = 17'b1010011001110011_0;
      patterns[3104] = 17'b1011011001110011_0;
      patterns[3105] = 17'b0101011001110000_0;
      patterns[3106] = 17'b0100011001110000_1;
      patterns[3107] = 17'b0000011000011100_0;
      patterns[3108] = 17'b1000011001110100_0;
      patterns[3109] = 17'b1001011001110100_0;
      patterns[3110] = 17'b1010011001110100_0;
      patterns[3111] = 17'b1011011001110100_0;
      patterns[3112] = 17'b0101011001110000_0;
      patterns[3113] = 17'b0100011001110000_1;
      patterns[3114] = 17'b0000011000001011_0;
      patterns[3115] = 17'b1000011001110101_0;
      patterns[3116] = 17'b1001011001110101_0;
      patterns[3117] = 17'b1010011001110101_0;
      patterns[3118] = 17'b1011011001110101_0;
      patterns[3119] = 17'b0101011001110000_0;
      patterns[3120] = 17'b0100011001110000_1;
      patterns[3121] = 17'b0000011011110100_0;
      patterns[3122] = 17'b1000011001110110_0;
      patterns[3123] = 17'b1001011001110110_0;
      patterns[3124] = 17'b1010011001110110_0;
      patterns[3125] = 17'b1011011001110110_0;
      patterns[3126] = 17'b0101011001110000_0;
      patterns[3127] = 17'b0100011001110000_1;
      patterns[3128] = 17'b0000011010111110_0;
      patterns[3129] = 17'b1000011001110111_0;
      patterns[3130] = 17'b1001011001110111_0;
      patterns[3131] = 17'b1010011001110111_0;
      patterns[3132] = 17'b1011011001110111_0;
      patterns[3133] = 17'b0101011001110000_0;
      patterns[3134] = 17'b0100011001110000_1;
      patterns[3135] = 17'b0000011000100101_0;
      patterns[3136] = 17'b1000011100000000_0;
      patterns[3137] = 17'b1001011100000000_0;
      patterns[3138] = 17'b1010011100000000_0;
      patterns[3139] = 17'b1011011100000000_0;
      patterns[3140] = 17'b0101011100000000_0;
      patterns[3141] = 17'b0100011100000000_1;
      patterns[3142] = 17'b0000011111111010_0;
      patterns[3143] = 17'b1000011100000001_0;
      patterns[3144] = 17'b1001011100000001_0;
      patterns[3145] = 17'b1010011100000001_0;
      patterns[3146] = 17'b1011011100000001_0;
      patterns[3147] = 17'b0101011100000000_0;
      patterns[3148] = 17'b0100011100000000_1;
      patterns[3149] = 17'b0000011101010000_0;
      patterns[3150] = 17'b1000011100000010_0;
      patterns[3151] = 17'b1001011100000010_0;
      patterns[3152] = 17'b1010011100000010_0;
      patterns[3153] = 17'b1011011100000010_0;
      patterns[3154] = 17'b0101011100000000_0;
      patterns[3155] = 17'b0100011100000000_1;
      patterns[3156] = 17'b0000011100100100_0;
      patterns[3157] = 17'b1000011100000011_0;
      patterns[3158] = 17'b1001011100000011_0;
      patterns[3159] = 17'b1010011100000011_0;
      patterns[3160] = 17'b1011011100000011_0;
      patterns[3161] = 17'b0101011100000000_0;
      patterns[3162] = 17'b0100011100000000_1;
      patterns[3163] = 17'b0000011111110010_0;
      patterns[3164] = 17'b1000011100000100_0;
      patterns[3165] = 17'b1001011100000100_0;
      patterns[3166] = 17'b1010011100000100_0;
      patterns[3167] = 17'b1011011100000100_0;
      patterns[3168] = 17'b0101011100000000_0;
      patterns[3169] = 17'b0100011100000000_1;
      patterns[3170] = 17'b0000011101011001_0;
      patterns[3171] = 17'b1000011100000101_0;
      patterns[3172] = 17'b1001011100000101_0;
      patterns[3173] = 17'b1010011100000101_0;
      patterns[3174] = 17'b1011011100000101_0;
      patterns[3175] = 17'b0101011100000000_0;
      patterns[3176] = 17'b0100011100000000_1;
      patterns[3177] = 17'b0000011100100100_0;
      patterns[3178] = 17'b1000011100000110_0;
      patterns[3179] = 17'b1001011100000110_0;
      patterns[3180] = 17'b1010011100000110_0;
      patterns[3181] = 17'b1011011100000110_0;
      patterns[3182] = 17'b0101011100000000_0;
      patterns[3183] = 17'b0100011100000000_1;
      patterns[3184] = 17'b0000011111110011_0;
      patterns[3185] = 17'b1000011100000111_0;
      patterns[3186] = 17'b1001011100000111_0;
      patterns[3187] = 17'b1010011100000111_0;
      patterns[3188] = 17'b1011011100000111_0;
      patterns[3189] = 17'b0101011100000000_0;
      patterns[3190] = 17'b0100011100000000_1;
      patterns[3191] = 17'b0000011100010110_0;
      patterns[3192] = 17'b1000011100010000_0;
      patterns[3193] = 17'b1001011100010000_0;
      patterns[3194] = 17'b1010011100010000_0;
      patterns[3195] = 17'b1011011100010000_0;
      patterns[3196] = 17'b0101011100010000_0;
      patterns[3197] = 17'b0100011100010000_1;
      patterns[3198] = 17'b0000011101100111_0;
      patterns[3199] = 17'b1000011100010001_0;
      patterns[3200] = 17'b1001011100010001_0;
      patterns[3201] = 17'b1010011100010001_0;
      patterns[3202] = 17'b1011011100010001_0;
      patterns[3203] = 17'b0101011100010000_0;
      patterns[3204] = 17'b0100011100010000_1;
      patterns[3205] = 17'b0000011111010100_0;
      patterns[3206] = 17'b1000011100010010_0;
      patterns[3207] = 17'b1001011100010010_0;
      patterns[3208] = 17'b1010011100010010_0;
      patterns[3209] = 17'b1011011100010010_0;
      patterns[3210] = 17'b0101011100010000_0;
      patterns[3211] = 17'b0100011100010000_1;
      patterns[3212] = 17'b0000011110100111_0;
      patterns[3213] = 17'b1000011100010011_0;
      patterns[3214] = 17'b1001011100010011_0;
      patterns[3215] = 17'b1010011100010011_0;
      patterns[3216] = 17'b1011011100010011_0;
      patterns[3217] = 17'b0101011100010000_0;
      patterns[3218] = 17'b0100011100010000_1;
      patterns[3219] = 17'b0000011101011001_0;
      patterns[3220] = 17'b1000011100010100_0;
      patterns[3221] = 17'b1001011100010100_0;
      patterns[3222] = 17'b1010011100010100_0;
      patterns[3223] = 17'b1011011100010100_0;
      patterns[3224] = 17'b0101011100010000_0;
      patterns[3225] = 17'b0100011100010000_1;
      patterns[3226] = 17'b0000011100100111_0;
      patterns[3227] = 17'b1000011100010101_0;
      patterns[3228] = 17'b1001011100010101_0;
      patterns[3229] = 17'b1010011100010101_0;
      patterns[3230] = 17'b1011011100010101_0;
      patterns[3231] = 17'b0101011100010000_0;
      patterns[3232] = 17'b0100011100010000_1;
      patterns[3233] = 17'b0000011110010001_0;
      patterns[3234] = 17'b1000011100010110_0;
      patterns[3235] = 17'b1001011100010110_0;
      patterns[3236] = 17'b1010011100010110_0;
      patterns[3237] = 17'b1011011100010110_0;
      patterns[3238] = 17'b0101011100010000_0;
      patterns[3239] = 17'b0100011100010000_1;
      patterns[3240] = 17'b0000011111010110_0;
      patterns[3241] = 17'b1000011100010111_0;
      patterns[3242] = 17'b1001011100010111_0;
      patterns[3243] = 17'b1010011100010111_0;
      patterns[3244] = 17'b1011011100010111_0;
      patterns[3245] = 17'b0101011100010000_0;
      patterns[3246] = 17'b0100011100010000_1;
      patterns[3247] = 17'b0000011110001011_0;
      patterns[3248] = 17'b1000011100100000_0;
      patterns[3249] = 17'b1001011100100000_0;
      patterns[3250] = 17'b1010011100100000_0;
      patterns[3251] = 17'b1011011100100000_0;
      patterns[3252] = 17'b0101011100100000_0;
      patterns[3253] = 17'b0100011100100000_1;
      patterns[3254] = 17'b0000011101101100_0;
      patterns[3255] = 17'b1000011100100001_0;
      patterns[3256] = 17'b1001011100100001_0;
      patterns[3257] = 17'b1010011100100001_0;
      patterns[3258] = 17'b1011011100100001_0;
      patterns[3259] = 17'b0101011100100000_0;
      patterns[3260] = 17'b0100011100100000_1;
      patterns[3261] = 17'b0000011101110100_0;
      patterns[3262] = 17'b1000011100100010_0;
      patterns[3263] = 17'b1001011100100010_0;
      patterns[3264] = 17'b1010011100100010_0;
      patterns[3265] = 17'b1011011100100010_0;
      patterns[3266] = 17'b0101011100100000_0;
      patterns[3267] = 17'b0100011100100000_1;
      patterns[3268] = 17'b0000011101110101_0;
      patterns[3269] = 17'b1000011100100011_0;
      patterns[3270] = 17'b1001011100100011_0;
      patterns[3271] = 17'b1010011100100011_0;
      patterns[3272] = 17'b1011011100100011_0;
      patterns[3273] = 17'b0101011100100000_0;
      patterns[3274] = 17'b0100011100100000_1;
      patterns[3275] = 17'b0000011110101100_0;
      patterns[3276] = 17'b1000011100100100_0;
      patterns[3277] = 17'b1001011100100100_0;
      patterns[3278] = 17'b1010011100100100_0;
      patterns[3279] = 17'b1011011100100100_0;
      patterns[3280] = 17'b0101011100100000_0;
      patterns[3281] = 17'b0100011100100000_1;
      patterns[3282] = 17'b0000011100011100_0;
      patterns[3283] = 17'b1000011100100101_0;
      patterns[3284] = 17'b1001011100100101_0;
      patterns[3285] = 17'b1010011100100101_0;
      patterns[3286] = 17'b1011011100100101_0;
      patterns[3287] = 17'b0101011100100000_0;
      patterns[3288] = 17'b0100011100100000_1;
      patterns[3289] = 17'b0000011110111101_0;
      patterns[3290] = 17'b1000011100100110_0;
      patterns[3291] = 17'b1001011100100110_0;
      patterns[3292] = 17'b1010011100100110_0;
      patterns[3293] = 17'b1011011100100110_0;
      patterns[3294] = 17'b0101011100100000_0;
      patterns[3295] = 17'b0100011100100000_1;
      patterns[3296] = 17'b0000011100001111_0;
      patterns[3297] = 17'b1000011100100111_0;
      patterns[3298] = 17'b1001011100100111_0;
      patterns[3299] = 17'b1010011100100111_0;
      patterns[3300] = 17'b1011011100100111_0;
      patterns[3301] = 17'b0101011100100000_0;
      patterns[3302] = 17'b0100011100100000_1;
      patterns[3303] = 17'b0000011110010010_0;
      patterns[3304] = 17'b1000011100110000_0;
      patterns[3305] = 17'b1001011100110000_0;
      patterns[3306] = 17'b1010011100110000_0;
      patterns[3307] = 17'b1011011100110000_0;
      patterns[3308] = 17'b0101011100110000_0;
      patterns[3309] = 17'b0100011100110000_1;
      patterns[3310] = 17'b0000011101110111_0;
      patterns[3311] = 17'b1000011100110001_0;
      patterns[3312] = 17'b1001011100110001_0;
      patterns[3313] = 17'b1010011100110001_0;
      patterns[3314] = 17'b1011011100110001_0;
      patterns[3315] = 17'b0101011100110000_0;
      patterns[3316] = 17'b0100011100110000_1;
      patterns[3317] = 17'b0000011101111111_0;
      patterns[3318] = 17'b1000011100110010_0;
      patterns[3319] = 17'b1001011100110010_0;
      patterns[3320] = 17'b1010011100110010_0;
      patterns[3321] = 17'b1011011100110010_0;
      patterns[3322] = 17'b0101011100110000_0;
      patterns[3323] = 17'b0100011100110000_1;
      patterns[3324] = 17'b0000011101101101_0;
      patterns[3325] = 17'b1000011100110011_0;
      patterns[3326] = 17'b1001011100110011_0;
      patterns[3327] = 17'b1010011100110011_0;
      patterns[3328] = 17'b1011011100110011_0;
      patterns[3329] = 17'b0101011100110000_0;
      patterns[3330] = 17'b0100011100110000_1;
      patterns[3331] = 17'b0000011100001010_0;
      patterns[3332] = 17'b1000011100110100_0;
      patterns[3333] = 17'b1001011100110100_0;
      patterns[3334] = 17'b1010011100110100_0;
      patterns[3335] = 17'b1011011100110100_0;
      patterns[3336] = 17'b0101011100110000_0;
      patterns[3337] = 17'b0100011100110000_1;
      patterns[3338] = 17'b0000011110100000_0;
      patterns[3339] = 17'b1000011100110101_0;
      patterns[3340] = 17'b1001011100110101_0;
      patterns[3341] = 17'b1010011100110101_0;
      patterns[3342] = 17'b1011011100110101_0;
      patterns[3343] = 17'b0101011100110000_0;
      patterns[3344] = 17'b0100011100110000_1;
      patterns[3345] = 17'b0000011100000000_0;
      patterns[3346] = 17'b1000011100110110_0;
      patterns[3347] = 17'b1001011100110110_0;
      patterns[3348] = 17'b1010011100110110_0;
      patterns[3349] = 17'b1011011100110110_0;
      patterns[3350] = 17'b0101011100110000_0;
      patterns[3351] = 17'b0100011100110000_1;
      patterns[3352] = 17'b0000011100010100_0;
      patterns[3353] = 17'b1000011100110111_0;
      patterns[3354] = 17'b1001011100110111_0;
      patterns[3355] = 17'b1010011100110111_0;
      patterns[3356] = 17'b1011011100110111_0;
      patterns[3357] = 17'b0101011100110000_0;
      patterns[3358] = 17'b0100011100110000_1;
      patterns[3359] = 17'b0000011110111100_0;
      patterns[3360] = 17'b1000011101000000_0;
      patterns[3361] = 17'b1001011101000000_0;
      patterns[3362] = 17'b1010011101000000_0;
      patterns[3363] = 17'b1011011101000000_0;
      patterns[3364] = 17'b0101011101000000_0;
      patterns[3365] = 17'b0100011101000000_1;
      patterns[3366] = 17'b0000011110111111_0;
      patterns[3367] = 17'b1000011101000001_0;
      patterns[3368] = 17'b1001011101000001_0;
      patterns[3369] = 17'b1010011101000001_0;
      patterns[3370] = 17'b1011011101000001_0;
      patterns[3371] = 17'b0101011101000000_0;
      patterns[3372] = 17'b0100011101000000_1;
      patterns[3373] = 17'b0000011100010011_0;
      patterns[3374] = 17'b1000011101000010_0;
      patterns[3375] = 17'b1001011101000010_0;
      patterns[3376] = 17'b1010011101000010_0;
      patterns[3377] = 17'b1011011101000010_0;
      patterns[3378] = 17'b0101011101000000_0;
      patterns[3379] = 17'b0100011101000000_1;
      patterns[3380] = 17'b0000011110011000_0;
      patterns[3381] = 17'b1000011101000011_0;
      patterns[3382] = 17'b1001011101000011_0;
      patterns[3383] = 17'b1010011101000011_0;
      patterns[3384] = 17'b1011011101000011_0;
      patterns[3385] = 17'b0101011101000000_0;
      patterns[3386] = 17'b0100011101000000_1;
      patterns[3387] = 17'b0000011100101001_0;
      patterns[3388] = 17'b1000011101000100_0;
      patterns[3389] = 17'b1001011101000100_0;
      patterns[3390] = 17'b1010011101000100_0;
      patterns[3391] = 17'b1011011101000100_0;
      patterns[3392] = 17'b0101011101000000_0;
      patterns[3393] = 17'b0100011101000000_1;
      patterns[3394] = 17'b0000011100010010_0;
      patterns[3395] = 17'b1000011101000101_0;
      patterns[3396] = 17'b1001011101000101_0;
      patterns[3397] = 17'b1010011101000101_0;
      patterns[3398] = 17'b1011011101000101_0;
      patterns[3399] = 17'b0101011101000000_0;
      patterns[3400] = 17'b0100011101000000_1;
      patterns[3401] = 17'b0000011111000110_0;
      patterns[3402] = 17'b1000011101000110_0;
      patterns[3403] = 17'b1001011101000110_0;
      patterns[3404] = 17'b1010011101000110_0;
      patterns[3405] = 17'b1011011101000110_0;
      patterns[3406] = 17'b0101011101000000_0;
      patterns[3407] = 17'b0100011101000000_1;
      patterns[3408] = 17'b0000011101100001_0;
      patterns[3409] = 17'b1000011101000111_0;
      patterns[3410] = 17'b1001011101000111_0;
      patterns[3411] = 17'b1010011101000111_0;
      patterns[3412] = 17'b1011011101000111_0;
      patterns[3413] = 17'b0101011101000000_0;
      patterns[3414] = 17'b0100011101000000_1;
      patterns[3415] = 17'b0000011101010011_0;
      patterns[3416] = 17'b1000011101010000_0;
      patterns[3417] = 17'b1001011101010000_0;
      patterns[3418] = 17'b1010011101010000_0;
      patterns[3419] = 17'b1011011101010000_0;
      patterns[3420] = 17'b0101011101010000_0;
      patterns[3421] = 17'b0100011101010000_1;
      patterns[3422] = 17'b0000011111101110_0;
      patterns[3423] = 17'b1000011101010001_0;
      patterns[3424] = 17'b1001011101010001_0;
      patterns[3425] = 17'b1010011101010001_0;
      patterns[3426] = 17'b1011011101010001_0;
      patterns[3427] = 17'b0101011101010000_0;
      patterns[3428] = 17'b0100011101010000_1;
      patterns[3429] = 17'b0000011111001000_0;
      patterns[3430] = 17'b1000011101010010_0;
      patterns[3431] = 17'b1001011101010010_0;
      patterns[3432] = 17'b1010011101010010_0;
      patterns[3433] = 17'b1011011101010010_0;
      patterns[3434] = 17'b0101011101010000_0;
      patterns[3435] = 17'b0100011101010000_1;
      patterns[3436] = 17'b0000011101111001_0;
      patterns[3437] = 17'b1000011101010011_0;
      patterns[3438] = 17'b1001011101010011_0;
      patterns[3439] = 17'b1010011101010011_0;
      patterns[3440] = 17'b1011011101010011_0;
      patterns[3441] = 17'b0101011101010000_0;
      patterns[3442] = 17'b0100011101010000_1;
      patterns[3443] = 17'b0000011111000100_0;
      patterns[3444] = 17'b1000011101010100_0;
      patterns[3445] = 17'b1001011101010100_0;
      patterns[3446] = 17'b1010011101010100_0;
      patterns[3447] = 17'b1011011101010100_0;
      patterns[3448] = 17'b0101011101010000_0;
      patterns[3449] = 17'b0100011101010000_1;
      patterns[3450] = 17'b0000011100110100_0;
      patterns[3451] = 17'b1000011101010101_0;
      patterns[3452] = 17'b1001011101010101_0;
      patterns[3453] = 17'b1010011101010101_0;
      patterns[3454] = 17'b1011011101010101_0;
      patterns[3455] = 17'b0101011101010000_0;
      patterns[3456] = 17'b0100011101010000_1;
      patterns[3457] = 17'b0000011111111100_0;
      patterns[3458] = 17'b1000011101010110_0;
      patterns[3459] = 17'b1001011101010110_0;
      patterns[3460] = 17'b1010011101010110_0;
      patterns[3461] = 17'b1011011101010110_0;
      patterns[3462] = 17'b0101011101010000_0;
      patterns[3463] = 17'b0100011101010000_1;
      patterns[3464] = 17'b0000011101001011_0;
      patterns[3465] = 17'b1000011101010111_0;
      patterns[3466] = 17'b1001011101010111_0;
      patterns[3467] = 17'b1010011101010111_0;
      patterns[3468] = 17'b1011011101010111_0;
      patterns[3469] = 17'b0101011101010000_0;
      patterns[3470] = 17'b0100011101010000_1;
      patterns[3471] = 17'b0000011100001110_0;
      patterns[3472] = 17'b1000011101100000_0;
      patterns[3473] = 17'b1001011101100000_0;
      patterns[3474] = 17'b1010011101100000_0;
      patterns[3475] = 17'b1011011101100000_0;
      patterns[3476] = 17'b0101011101100000_0;
      patterns[3477] = 17'b0100011101100000_1;
      patterns[3478] = 17'b0000011100010100_0;
      patterns[3479] = 17'b1000011101100001_0;
      patterns[3480] = 17'b1001011101100001_0;
      patterns[3481] = 17'b1010011101100001_0;
      patterns[3482] = 17'b1011011101100001_0;
      patterns[3483] = 17'b0101011101100000_0;
      patterns[3484] = 17'b0100011101100000_1;
      patterns[3485] = 17'b0000011111110101_0;
      patterns[3486] = 17'b1000011101100010_0;
      patterns[3487] = 17'b1001011101100010_0;
      patterns[3488] = 17'b1010011101100010_0;
      patterns[3489] = 17'b1011011101100010_0;
      patterns[3490] = 17'b0101011101100000_0;
      patterns[3491] = 17'b0100011101100000_1;
      patterns[3492] = 17'b0000011111001001_0;
      patterns[3493] = 17'b1000011101100011_0;
      patterns[3494] = 17'b1001011101100011_0;
      patterns[3495] = 17'b1010011101100011_0;
      patterns[3496] = 17'b1011011101100011_0;
      patterns[3497] = 17'b0101011101100000_0;
      patterns[3498] = 17'b0100011101100000_1;
      patterns[3499] = 17'b0000011111101000_0;
      patterns[3500] = 17'b1000011101100100_0;
      patterns[3501] = 17'b1001011101100100_0;
      patterns[3502] = 17'b1010011101100100_0;
      patterns[3503] = 17'b1011011101100100_0;
      patterns[3504] = 17'b0101011101100000_0;
      patterns[3505] = 17'b0100011101100000_1;
      patterns[3506] = 17'b0000011111110010_0;
      patterns[3507] = 17'b1000011101100101_0;
      patterns[3508] = 17'b1001011101100101_0;
      patterns[3509] = 17'b1010011101100101_0;
      patterns[3510] = 17'b1011011101100101_0;
      patterns[3511] = 17'b0101011101100000_0;
      patterns[3512] = 17'b0100011101100000_1;
      patterns[3513] = 17'b0000011100001001_0;
      patterns[3514] = 17'b1000011101100110_0;
      patterns[3515] = 17'b1001011101100110_0;
      patterns[3516] = 17'b1010011101100110_0;
      patterns[3517] = 17'b1011011101100110_0;
      patterns[3518] = 17'b0101011101100000_0;
      patterns[3519] = 17'b0100011101100000_1;
      patterns[3520] = 17'b0000011100100101_0;
      patterns[3521] = 17'b1000011101100111_0;
      patterns[3522] = 17'b1001011101100111_0;
      patterns[3523] = 17'b1010011101100111_0;
      patterns[3524] = 17'b1011011101100111_0;
      patterns[3525] = 17'b0101011101100000_0;
      patterns[3526] = 17'b0100011101100000_1;
      patterns[3527] = 17'b0000011110100010_0;
      patterns[3528] = 17'b1000011101110000_0;
      patterns[3529] = 17'b1001011101110000_0;
      patterns[3530] = 17'b1010011101110000_0;
      patterns[3531] = 17'b1011011101110000_0;
      patterns[3532] = 17'b0101011101110000_0;
      patterns[3533] = 17'b0100011101110000_1;
      patterns[3534] = 17'b0000011100101001_0;
      patterns[3535] = 17'b1000011101110001_0;
      patterns[3536] = 17'b1001011101110001_0;
      patterns[3537] = 17'b1010011101110001_0;
      patterns[3538] = 17'b1011011101110001_0;
      patterns[3539] = 17'b0101011101110000_0;
      patterns[3540] = 17'b0100011101110000_1;
      patterns[3541] = 17'b0000011100010011_0;
      patterns[3542] = 17'b1000011101110010_0;
      patterns[3543] = 17'b1001011101110010_0;
      patterns[3544] = 17'b1010011101110010_0;
      patterns[3545] = 17'b1011011101110010_0;
      patterns[3546] = 17'b0101011101110000_0;
      patterns[3547] = 17'b0100011101110000_1;
      patterns[3548] = 17'b0000011110010011_0;
      patterns[3549] = 17'b1000011101110011_0;
      patterns[3550] = 17'b1001011101110011_0;
      patterns[3551] = 17'b1010011101110011_0;
      patterns[3552] = 17'b1011011101110011_0;
      patterns[3553] = 17'b0101011101110000_0;
      patterns[3554] = 17'b0100011101110000_1;
      patterns[3555] = 17'b0000011110111011_0;
      patterns[3556] = 17'b1000011101110100_0;
      patterns[3557] = 17'b1001011101110100_0;
      patterns[3558] = 17'b1010011101110100_0;
      patterns[3559] = 17'b1011011101110100_0;
      patterns[3560] = 17'b0101011101110000_0;
      patterns[3561] = 17'b0100011101110000_1;
      patterns[3562] = 17'b0000011100001010_0;
      patterns[3563] = 17'b1000011101110101_0;
      patterns[3564] = 17'b1001011101110101_0;
      patterns[3565] = 17'b1010011101110101_0;
      patterns[3566] = 17'b1011011101110101_0;
      patterns[3567] = 17'b0101011101110000_0;
      patterns[3568] = 17'b0100011101110000_1;
      patterns[3569] = 17'b0000011100001011_0;
      patterns[3570] = 17'b1000011101110110_0;
      patterns[3571] = 17'b1001011101110110_0;
      patterns[3572] = 17'b1010011101110110_0;
      patterns[3573] = 17'b1011011101110110_0;
      patterns[3574] = 17'b0101011101110000_0;
      patterns[3575] = 17'b0100011101110000_1;
      patterns[3576] = 17'b0000011111001111_0;
      patterns[3577] = 17'b1000011101110111_0;
      patterns[3578] = 17'b1001011101110111_0;
      patterns[3579] = 17'b1010011101110111_0;
      patterns[3580] = 17'b1011011101110111_0;
      patterns[3581] = 17'b0101011101110000_0;
      patterns[3582] = 17'b0100011101110000_1;
      patterns[3583] = 17'b0000011111110100_0;

      for (i = 0; i < 3584; i = i + 1)
      begin
        INST = patterns[i][16:1];
        #10;
        if (patterns[i][0] !== 1'hx)
        begin
          if (STR !== patterns[i][0])
          begin
            $display("%d:STR: (assertion error). Expected %h, found %h", i, patterns[i][0], STR);
            $finish;
          end
        end
      end

      $display("All tests passed.");
    end
    endmodule
