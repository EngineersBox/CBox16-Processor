//  A testbench for control_unit_ALUOP_tb
`timescale 1us/1ns

module control_unit_ALUOP_tb;
    reg [15:0] INST;
    reg FL_Z;
    wire [1:0] ALUOP;
    wire [2:0] RS1;
    wire [2:0] RS2;
    wire [2:0] WS;
    wire STR;
    wire WE;
    wire [1:0] DMUX;
    wire LDR;
    wire FL_EN;
    wire HE;

  control_unit control_unit0 (
    .INST(INST),
    .FL_Z(FL_Z),
    .ALUOP(ALUOP),
    .RS1(RS1),
    .RS2(RS2),
    .WS(WS),
    .STR(STR),
    .WE(WE),
    .DMUX(DMUX),
    .LDR(LDR),
    .FL_EN(FL_EN),
    .HE(HE)
  );

    reg [17:0] patterns[0:2047];
    integer i;

    initial begin
      patterns[0] = 18'b1000000000000000_00;
      patterns[1] = 18'b1001000000000000_01;
      patterns[2] = 18'b1010000000000000_10;
      patterns[3] = 18'b1011000000000000_11;
      patterns[4] = 18'b1000000000000001_00;
      patterns[5] = 18'b1001000000000001_01;
      patterns[6] = 18'b1010000000000001_10;
      patterns[7] = 18'b1011000000000001_11;
      patterns[8] = 18'b1000000000000010_00;
      patterns[9] = 18'b1001000000000010_01;
      patterns[10] = 18'b1010000000000010_10;
      patterns[11] = 18'b1011000000000010_11;
      patterns[12] = 18'b1000000000000011_00;
      patterns[13] = 18'b1001000000000011_01;
      patterns[14] = 18'b1010000000000011_10;
      patterns[15] = 18'b1011000000000011_11;
      patterns[16] = 18'b1000000000000100_00;
      patterns[17] = 18'b1001000000000100_01;
      patterns[18] = 18'b1010000000000100_10;
      patterns[19] = 18'b1011000000000100_11;
      patterns[20] = 18'b1000000000000101_00;
      patterns[21] = 18'b1001000000000101_01;
      patterns[22] = 18'b1010000000000101_10;
      patterns[23] = 18'b1011000000000101_11;
      patterns[24] = 18'b1000000000000110_00;
      patterns[25] = 18'b1001000000000110_01;
      patterns[26] = 18'b1010000000000110_10;
      patterns[27] = 18'b1011000000000110_11;
      patterns[28] = 18'b1000000000000111_00;
      patterns[29] = 18'b1001000000000111_01;
      patterns[30] = 18'b1010000000000111_10;
      patterns[31] = 18'b1011000000000111_11;
      patterns[32] = 18'b1000000000010000_00;
      patterns[33] = 18'b1001000000010000_01;
      patterns[34] = 18'b1010000000010000_10;
      patterns[35] = 18'b1011000000010000_11;
      patterns[36] = 18'b1000000000010001_00;
      patterns[37] = 18'b1001000000010001_01;
      patterns[38] = 18'b1010000000010001_10;
      patterns[39] = 18'b1011000000010001_11;
      patterns[40] = 18'b1000000000010010_00;
      patterns[41] = 18'b1001000000010010_01;
      patterns[42] = 18'b1010000000010010_10;
      patterns[43] = 18'b1011000000010010_11;
      patterns[44] = 18'b1000000000010011_00;
      patterns[45] = 18'b1001000000010011_01;
      patterns[46] = 18'b1010000000010011_10;
      patterns[47] = 18'b1011000000010011_11;
      patterns[48] = 18'b1000000000010100_00;
      patterns[49] = 18'b1001000000010100_01;
      patterns[50] = 18'b1010000000010100_10;
      patterns[51] = 18'b1011000000010100_11;
      patterns[52] = 18'b1000000000010101_00;
      patterns[53] = 18'b1001000000010101_01;
      patterns[54] = 18'b1010000000010101_10;
      patterns[55] = 18'b1011000000010101_11;
      patterns[56] = 18'b1000000000010110_00;
      patterns[57] = 18'b1001000000010110_01;
      patterns[58] = 18'b1010000000010110_10;
      patterns[59] = 18'b1011000000010110_11;
      patterns[60] = 18'b1000000000010111_00;
      patterns[61] = 18'b1001000000010111_01;
      patterns[62] = 18'b1010000000010111_10;
      patterns[63] = 18'b1011000000010111_11;
      patterns[64] = 18'b1000000000100000_00;
      patterns[65] = 18'b1001000000100000_01;
      patterns[66] = 18'b1010000000100000_10;
      patterns[67] = 18'b1011000000100000_11;
      patterns[68] = 18'b1000000000100001_00;
      patterns[69] = 18'b1001000000100001_01;
      patterns[70] = 18'b1010000000100001_10;
      patterns[71] = 18'b1011000000100001_11;
      patterns[72] = 18'b1000000000100010_00;
      patterns[73] = 18'b1001000000100010_01;
      patterns[74] = 18'b1010000000100010_10;
      patterns[75] = 18'b1011000000100010_11;
      patterns[76] = 18'b1000000000100011_00;
      patterns[77] = 18'b1001000000100011_01;
      patterns[78] = 18'b1010000000100011_10;
      patterns[79] = 18'b1011000000100011_11;
      patterns[80] = 18'b1000000000100100_00;
      patterns[81] = 18'b1001000000100100_01;
      patterns[82] = 18'b1010000000100100_10;
      patterns[83] = 18'b1011000000100100_11;
      patterns[84] = 18'b1000000000100101_00;
      patterns[85] = 18'b1001000000100101_01;
      patterns[86] = 18'b1010000000100101_10;
      patterns[87] = 18'b1011000000100101_11;
      patterns[88] = 18'b1000000000100110_00;
      patterns[89] = 18'b1001000000100110_01;
      patterns[90] = 18'b1010000000100110_10;
      patterns[91] = 18'b1011000000100110_11;
      patterns[92] = 18'b1000000000100111_00;
      patterns[93] = 18'b1001000000100111_01;
      patterns[94] = 18'b1010000000100111_10;
      patterns[95] = 18'b1011000000100111_11;
      patterns[96] = 18'b1000000000110000_00;
      patterns[97] = 18'b1001000000110000_01;
      patterns[98] = 18'b1010000000110000_10;
      patterns[99] = 18'b1011000000110000_11;
      patterns[100] = 18'b1000000000110001_00;
      patterns[101] = 18'b1001000000110001_01;
      patterns[102] = 18'b1010000000110001_10;
      patterns[103] = 18'b1011000000110001_11;
      patterns[104] = 18'b1000000000110010_00;
      patterns[105] = 18'b1001000000110010_01;
      patterns[106] = 18'b1010000000110010_10;
      patterns[107] = 18'b1011000000110010_11;
      patterns[108] = 18'b1000000000110011_00;
      patterns[109] = 18'b1001000000110011_01;
      patterns[110] = 18'b1010000000110011_10;
      patterns[111] = 18'b1011000000110011_11;
      patterns[112] = 18'b1000000000110100_00;
      patterns[113] = 18'b1001000000110100_01;
      patterns[114] = 18'b1010000000110100_10;
      patterns[115] = 18'b1011000000110100_11;
      patterns[116] = 18'b1000000000110101_00;
      patterns[117] = 18'b1001000000110101_01;
      patterns[118] = 18'b1010000000110101_10;
      patterns[119] = 18'b1011000000110101_11;
      patterns[120] = 18'b1000000000110110_00;
      patterns[121] = 18'b1001000000110110_01;
      patterns[122] = 18'b1010000000110110_10;
      patterns[123] = 18'b1011000000110110_11;
      patterns[124] = 18'b1000000000110111_00;
      patterns[125] = 18'b1001000000110111_01;
      patterns[126] = 18'b1010000000110111_10;
      patterns[127] = 18'b1011000000110111_11;
      patterns[128] = 18'b1000000001000000_00;
      patterns[129] = 18'b1001000001000000_01;
      patterns[130] = 18'b1010000001000000_10;
      patterns[131] = 18'b1011000001000000_11;
      patterns[132] = 18'b1000000001000001_00;
      patterns[133] = 18'b1001000001000001_01;
      patterns[134] = 18'b1010000001000001_10;
      patterns[135] = 18'b1011000001000001_11;
      patterns[136] = 18'b1000000001000010_00;
      patterns[137] = 18'b1001000001000010_01;
      patterns[138] = 18'b1010000001000010_10;
      patterns[139] = 18'b1011000001000010_11;
      patterns[140] = 18'b1000000001000011_00;
      patterns[141] = 18'b1001000001000011_01;
      patterns[142] = 18'b1010000001000011_10;
      patterns[143] = 18'b1011000001000011_11;
      patterns[144] = 18'b1000000001000100_00;
      patterns[145] = 18'b1001000001000100_01;
      patterns[146] = 18'b1010000001000100_10;
      patterns[147] = 18'b1011000001000100_11;
      patterns[148] = 18'b1000000001000101_00;
      patterns[149] = 18'b1001000001000101_01;
      patterns[150] = 18'b1010000001000101_10;
      patterns[151] = 18'b1011000001000101_11;
      patterns[152] = 18'b1000000001000110_00;
      patterns[153] = 18'b1001000001000110_01;
      patterns[154] = 18'b1010000001000110_10;
      patterns[155] = 18'b1011000001000110_11;
      patterns[156] = 18'b1000000001000111_00;
      patterns[157] = 18'b1001000001000111_01;
      patterns[158] = 18'b1010000001000111_10;
      patterns[159] = 18'b1011000001000111_11;
      patterns[160] = 18'b1000000001010000_00;
      patterns[161] = 18'b1001000001010000_01;
      patterns[162] = 18'b1010000001010000_10;
      patterns[163] = 18'b1011000001010000_11;
      patterns[164] = 18'b1000000001010001_00;
      patterns[165] = 18'b1001000001010001_01;
      patterns[166] = 18'b1010000001010001_10;
      patterns[167] = 18'b1011000001010001_11;
      patterns[168] = 18'b1000000001010010_00;
      patterns[169] = 18'b1001000001010010_01;
      patterns[170] = 18'b1010000001010010_10;
      patterns[171] = 18'b1011000001010010_11;
      patterns[172] = 18'b1000000001010011_00;
      patterns[173] = 18'b1001000001010011_01;
      patterns[174] = 18'b1010000001010011_10;
      patterns[175] = 18'b1011000001010011_11;
      patterns[176] = 18'b1000000001010100_00;
      patterns[177] = 18'b1001000001010100_01;
      patterns[178] = 18'b1010000001010100_10;
      patterns[179] = 18'b1011000001010100_11;
      patterns[180] = 18'b1000000001010101_00;
      patterns[181] = 18'b1001000001010101_01;
      patterns[182] = 18'b1010000001010101_10;
      patterns[183] = 18'b1011000001010101_11;
      patterns[184] = 18'b1000000001010110_00;
      patterns[185] = 18'b1001000001010110_01;
      patterns[186] = 18'b1010000001010110_10;
      patterns[187] = 18'b1011000001010110_11;
      patterns[188] = 18'b1000000001010111_00;
      patterns[189] = 18'b1001000001010111_01;
      patterns[190] = 18'b1010000001010111_10;
      patterns[191] = 18'b1011000001010111_11;
      patterns[192] = 18'b1000000001100000_00;
      patterns[193] = 18'b1001000001100000_01;
      patterns[194] = 18'b1010000001100000_10;
      patterns[195] = 18'b1011000001100000_11;
      patterns[196] = 18'b1000000001100001_00;
      patterns[197] = 18'b1001000001100001_01;
      patterns[198] = 18'b1010000001100001_10;
      patterns[199] = 18'b1011000001100001_11;
      patterns[200] = 18'b1000000001100010_00;
      patterns[201] = 18'b1001000001100010_01;
      patterns[202] = 18'b1010000001100010_10;
      patterns[203] = 18'b1011000001100010_11;
      patterns[204] = 18'b1000000001100011_00;
      patterns[205] = 18'b1001000001100011_01;
      patterns[206] = 18'b1010000001100011_10;
      patterns[207] = 18'b1011000001100011_11;
      patterns[208] = 18'b1000000001100100_00;
      patterns[209] = 18'b1001000001100100_01;
      patterns[210] = 18'b1010000001100100_10;
      patterns[211] = 18'b1011000001100100_11;
      patterns[212] = 18'b1000000001100101_00;
      patterns[213] = 18'b1001000001100101_01;
      patterns[214] = 18'b1010000001100101_10;
      patterns[215] = 18'b1011000001100101_11;
      patterns[216] = 18'b1000000001100110_00;
      patterns[217] = 18'b1001000001100110_01;
      patterns[218] = 18'b1010000001100110_10;
      patterns[219] = 18'b1011000001100110_11;
      patterns[220] = 18'b1000000001100111_00;
      patterns[221] = 18'b1001000001100111_01;
      patterns[222] = 18'b1010000001100111_10;
      patterns[223] = 18'b1011000001100111_11;
      patterns[224] = 18'b1000000001110000_00;
      patterns[225] = 18'b1001000001110000_01;
      patterns[226] = 18'b1010000001110000_10;
      patterns[227] = 18'b1011000001110000_11;
      patterns[228] = 18'b1000000001110001_00;
      patterns[229] = 18'b1001000001110001_01;
      patterns[230] = 18'b1010000001110001_10;
      patterns[231] = 18'b1011000001110001_11;
      patterns[232] = 18'b1000000001110010_00;
      patterns[233] = 18'b1001000001110010_01;
      patterns[234] = 18'b1010000001110010_10;
      patterns[235] = 18'b1011000001110010_11;
      patterns[236] = 18'b1000000001110011_00;
      patterns[237] = 18'b1001000001110011_01;
      patterns[238] = 18'b1010000001110011_10;
      patterns[239] = 18'b1011000001110011_11;
      patterns[240] = 18'b1000000001110100_00;
      patterns[241] = 18'b1001000001110100_01;
      patterns[242] = 18'b1010000001110100_10;
      patterns[243] = 18'b1011000001110100_11;
      patterns[244] = 18'b1000000001110101_00;
      patterns[245] = 18'b1001000001110101_01;
      patterns[246] = 18'b1010000001110101_10;
      patterns[247] = 18'b1011000001110101_11;
      patterns[248] = 18'b1000000001110110_00;
      patterns[249] = 18'b1001000001110110_01;
      patterns[250] = 18'b1010000001110110_10;
      patterns[251] = 18'b1011000001110110_11;
      patterns[252] = 18'b1000000001110111_00;
      patterns[253] = 18'b1001000001110111_01;
      patterns[254] = 18'b1010000001110111_10;
      patterns[255] = 18'b1011000001110111_11;
      patterns[256] = 18'b1000000100000000_00;
      patterns[257] = 18'b1001000100000000_01;
      patterns[258] = 18'b1010000100000000_10;
      patterns[259] = 18'b1011000100000000_11;
      patterns[260] = 18'b1000000100000001_00;
      patterns[261] = 18'b1001000100000001_01;
      patterns[262] = 18'b1010000100000001_10;
      patterns[263] = 18'b1011000100000001_11;
      patterns[264] = 18'b1000000100000010_00;
      patterns[265] = 18'b1001000100000010_01;
      patterns[266] = 18'b1010000100000010_10;
      patterns[267] = 18'b1011000100000010_11;
      patterns[268] = 18'b1000000100000011_00;
      patterns[269] = 18'b1001000100000011_01;
      patterns[270] = 18'b1010000100000011_10;
      patterns[271] = 18'b1011000100000011_11;
      patterns[272] = 18'b1000000100000100_00;
      patterns[273] = 18'b1001000100000100_01;
      patterns[274] = 18'b1010000100000100_10;
      patterns[275] = 18'b1011000100000100_11;
      patterns[276] = 18'b1000000100000101_00;
      patterns[277] = 18'b1001000100000101_01;
      patterns[278] = 18'b1010000100000101_10;
      patterns[279] = 18'b1011000100000101_11;
      patterns[280] = 18'b1000000100000110_00;
      patterns[281] = 18'b1001000100000110_01;
      patterns[282] = 18'b1010000100000110_10;
      patterns[283] = 18'b1011000100000110_11;
      patterns[284] = 18'b1000000100000111_00;
      patterns[285] = 18'b1001000100000111_01;
      patterns[286] = 18'b1010000100000111_10;
      patterns[287] = 18'b1011000100000111_11;
      patterns[288] = 18'b1000000100010000_00;
      patterns[289] = 18'b1001000100010000_01;
      patterns[290] = 18'b1010000100010000_10;
      patterns[291] = 18'b1011000100010000_11;
      patterns[292] = 18'b1000000100010001_00;
      patterns[293] = 18'b1001000100010001_01;
      patterns[294] = 18'b1010000100010001_10;
      patterns[295] = 18'b1011000100010001_11;
      patterns[296] = 18'b1000000100010010_00;
      patterns[297] = 18'b1001000100010010_01;
      patterns[298] = 18'b1010000100010010_10;
      patterns[299] = 18'b1011000100010010_11;
      patterns[300] = 18'b1000000100010011_00;
      patterns[301] = 18'b1001000100010011_01;
      patterns[302] = 18'b1010000100010011_10;
      patterns[303] = 18'b1011000100010011_11;
      patterns[304] = 18'b1000000100010100_00;
      patterns[305] = 18'b1001000100010100_01;
      patterns[306] = 18'b1010000100010100_10;
      patterns[307] = 18'b1011000100010100_11;
      patterns[308] = 18'b1000000100010101_00;
      patterns[309] = 18'b1001000100010101_01;
      patterns[310] = 18'b1010000100010101_10;
      patterns[311] = 18'b1011000100010101_11;
      patterns[312] = 18'b1000000100010110_00;
      patterns[313] = 18'b1001000100010110_01;
      patterns[314] = 18'b1010000100010110_10;
      patterns[315] = 18'b1011000100010110_11;
      patterns[316] = 18'b1000000100010111_00;
      patterns[317] = 18'b1001000100010111_01;
      patterns[318] = 18'b1010000100010111_10;
      patterns[319] = 18'b1011000100010111_11;
      patterns[320] = 18'b1000000100100000_00;
      patterns[321] = 18'b1001000100100000_01;
      patterns[322] = 18'b1010000100100000_10;
      patterns[323] = 18'b1011000100100000_11;
      patterns[324] = 18'b1000000100100001_00;
      patterns[325] = 18'b1001000100100001_01;
      patterns[326] = 18'b1010000100100001_10;
      patterns[327] = 18'b1011000100100001_11;
      patterns[328] = 18'b1000000100100010_00;
      patterns[329] = 18'b1001000100100010_01;
      patterns[330] = 18'b1010000100100010_10;
      patterns[331] = 18'b1011000100100010_11;
      patterns[332] = 18'b1000000100100011_00;
      patterns[333] = 18'b1001000100100011_01;
      patterns[334] = 18'b1010000100100011_10;
      patterns[335] = 18'b1011000100100011_11;
      patterns[336] = 18'b1000000100100100_00;
      patterns[337] = 18'b1001000100100100_01;
      patterns[338] = 18'b1010000100100100_10;
      patterns[339] = 18'b1011000100100100_11;
      patterns[340] = 18'b1000000100100101_00;
      patterns[341] = 18'b1001000100100101_01;
      patterns[342] = 18'b1010000100100101_10;
      patterns[343] = 18'b1011000100100101_11;
      patterns[344] = 18'b1000000100100110_00;
      patterns[345] = 18'b1001000100100110_01;
      patterns[346] = 18'b1010000100100110_10;
      patterns[347] = 18'b1011000100100110_11;
      patterns[348] = 18'b1000000100100111_00;
      patterns[349] = 18'b1001000100100111_01;
      patterns[350] = 18'b1010000100100111_10;
      patterns[351] = 18'b1011000100100111_11;
      patterns[352] = 18'b1000000100110000_00;
      patterns[353] = 18'b1001000100110000_01;
      patterns[354] = 18'b1010000100110000_10;
      patterns[355] = 18'b1011000100110000_11;
      patterns[356] = 18'b1000000100110001_00;
      patterns[357] = 18'b1001000100110001_01;
      patterns[358] = 18'b1010000100110001_10;
      patterns[359] = 18'b1011000100110001_11;
      patterns[360] = 18'b1000000100110010_00;
      patterns[361] = 18'b1001000100110010_01;
      patterns[362] = 18'b1010000100110010_10;
      patterns[363] = 18'b1011000100110010_11;
      patterns[364] = 18'b1000000100110011_00;
      patterns[365] = 18'b1001000100110011_01;
      patterns[366] = 18'b1010000100110011_10;
      patterns[367] = 18'b1011000100110011_11;
      patterns[368] = 18'b1000000100110100_00;
      patterns[369] = 18'b1001000100110100_01;
      patterns[370] = 18'b1010000100110100_10;
      patterns[371] = 18'b1011000100110100_11;
      patterns[372] = 18'b1000000100110101_00;
      patterns[373] = 18'b1001000100110101_01;
      patterns[374] = 18'b1010000100110101_10;
      patterns[375] = 18'b1011000100110101_11;
      patterns[376] = 18'b1000000100110110_00;
      patterns[377] = 18'b1001000100110110_01;
      patterns[378] = 18'b1010000100110110_10;
      patterns[379] = 18'b1011000100110110_11;
      patterns[380] = 18'b1000000100110111_00;
      patterns[381] = 18'b1001000100110111_01;
      patterns[382] = 18'b1010000100110111_10;
      patterns[383] = 18'b1011000100110111_11;
      patterns[384] = 18'b1000000101000000_00;
      patterns[385] = 18'b1001000101000000_01;
      patterns[386] = 18'b1010000101000000_10;
      patterns[387] = 18'b1011000101000000_11;
      patterns[388] = 18'b1000000101000001_00;
      patterns[389] = 18'b1001000101000001_01;
      patterns[390] = 18'b1010000101000001_10;
      patterns[391] = 18'b1011000101000001_11;
      patterns[392] = 18'b1000000101000010_00;
      patterns[393] = 18'b1001000101000010_01;
      patterns[394] = 18'b1010000101000010_10;
      patterns[395] = 18'b1011000101000010_11;
      patterns[396] = 18'b1000000101000011_00;
      patterns[397] = 18'b1001000101000011_01;
      patterns[398] = 18'b1010000101000011_10;
      patterns[399] = 18'b1011000101000011_11;
      patterns[400] = 18'b1000000101000100_00;
      patterns[401] = 18'b1001000101000100_01;
      patterns[402] = 18'b1010000101000100_10;
      patterns[403] = 18'b1011000101000100_11;
      patterns[404] = 18'b1000000101000101_00;
      patterns[405] = 18'b1001000101000101_01;
      patterns[406] = 18'b1010000101000101_10;
      patterns[407] = 18'b1011000101000101_11;
      patterns[408] = 18'b1000000101000110_00;
      patterns[409] = 18'b1001000101000110_01;
      patterns[410] = 18'b1010000101000110_10;
      patterns[411] = 18'b1011000101000110_11;
      patterns[412] = 18'b1000000101000111_00;
      patterns[413] = 18'b1001000101000111_01;
      patterns[414] = 18'b1010000101000111_10;
      patterns[415] = 18'b1011000101000111_11;
      patterns[416] = 18'b1000000101010000_00;
      patterns[417] = 18'b1001000101010000_01;
      patterns[418] = 18'b1010000101010000_10;
      patterns[419] = 18'b1011000101010000_11;
      patterns[420] = 18'b1000000101010001_00;
      patterns[421] = 18'b1001000101010001_01;
      patterns[422] = 18'b1010000101010001_10;
      patterns[423] = 18'b1011000101010001_11;
      patterns[424] = 18'b1000000101010010_00;
      patterns[425] = 18'b1001000101010010_01;
      patterns[426] = 18'b1010000101010010_10;
      patterns[427] = 18'b1011000101010010_11;
      patterns[428] = 18'b1000000101010011_00;
      patterns[429] = 18'b1001000101010011_01;
      patterns[430] = 18'b1010000101010011_10;
      patterns[431] = 18'b1011000101010011_11;
      patterns[432] = 18'b1000000101010100_00;
      patterns[433] = 18'b1001000101010100_01;
      patterns[434] = 18'b1010000101010100_10;
      patterns[435] = 18'b1011000101010100_11;
      patterns[436] = 18'b1000000101010101_00;
      patterns[437] = 18'b1001000101010101_01;
      patterns[438] = 18'b1010000101010101_10;
      patterns[439] = 18'b1011000101010101_11;
      patterns[440] = 18'b1000000101010110_00;
      patterns[441] = 18'b1001000101010110_01;
      patterns[442] = 18'b1010000101010110_10;
      patterns[443] = 18'b1011000101010110_11;
      patterns[444] = 18'b1000000101010111_00;
      patterns[445] = 18'b1001000101010111_01;
      patterns[446] = 18'b1010000101010111_10;
      patterns[447] = 18'b1011000101010111_11;
      patterns[448] = 18'b1000000101100000_00;
      patterns[449] = 18'b1001000101100000_01;
      patterns[450] = 18'b1010000101100000_10;
      patterns[451] = 18'b1011000101100000_11;
      patterns[452] = 18'b1000000101100001_00;
      patterns[453] = 18'b1001000101100001_01;
      patterns[454] = 18'b1010000101100001_10;
      patterns[455] = 18'b1011000101100001_11;
      patterns[456] = 18'b1000000101100010_00;
      patterns[457] = 18'b1001000101100010_01;
      patterns[458] = 18'b1010000101100010_10;
      patterns[459] = 18'b1011000101100010_11;
      patterns[460] = 18'b1000000101100011_00;
      patterns[461] = 18'b1001000101100011_01;
      patterns[462] = 18'b1010000101100011_10;
      patterns[463] = 18'b1011000101100011_11;
      patterns[464] = 18'b1000000101100100_00;
      patterns[465] = 18'b1001000101100100_01;
      patterns[466] = 18'b1010000101100100_10;
      patterns[467] = 18'b1011000101100100_11;
      patterns[468] = 18'b1000000101100101_00;
      patterns[469] = 18'b1001000101100101_01;
      patterns[470] = 18'b1010000101100101_10;
      patterns[471] = 18'b1011000101100101_11;
      patterns[472] = 18'b1000000101100110_00;
      patterns[473] = 18'b1001000101100110_01;
      patterns[474] = 18'b1010000101100110_10;
      patterns[475] = 18'b1011000101100110_11;
      patterns[476] = 18'b1000000101100111_00;
      patterns[477] = 18'b1001000101100111_01;
      patterns[478] = 18'b1010000101100111_10;
      patterns[479] = 18'b1011000101100111_11;
      patterns[480] = 18'b1000000101110000_00;
      patterns[481] = 18'b1001000101110000_01;
      patterns[482] = 18'b1010000101110000_10;
      patterns[483] = 18'b1011000101110000_11;
      patterns[484] = 18'b1000000101110001_00;
      patterns[485] = 18'b1001000101110001_01;
      patterns[486] = 18'b1010000101110001_10;
      patterns[487] = 18'b1011000101110001_11;
      patterns[488] = 18'b1000000101110010_00;
      patterns[489] = 18'b1001000101110010_01;
      patterns[490] = 18'b1010000101110010_10;
      patterns[491] = 18'b1011000101110010_11;
      patterns[492] = 18'b1000000101110011_00;
      patterns[493] = 18'b1001000101110011_01;
      patterns[494] = 18'b1010000101110011_10;
      patterns[495] = 18'b1011000101110011_11;
      patterns[496] = 18'b1000000101110100_00;
      patterns[497] = 18'b1001000101110100_01;
      patterns[498] = 18'b1010000101110100_10;
      patterns[499] = 18'b1011000101110100_11;
      patterns[500] = 18'b1000000101110101_00;
      patterns[501] = 18'b1001000101110101_01;
      patterns[502] = 18'b1010000101110101_10;
      patterns[503] = 18'b1011000101110101_11;
      patterns[504] = 18'b1000000101110110_00;
      patterns[505] = 18'b1001000101110110_01;
      patterns[506] = 18'b1010000101110110_10;
      patterns[507] = 18'b1011000101110110_11;
      patterns[508] = 18'b1000000101110111_00;
      patterns[509] = 18'b1001000101110111_01;
      patterns[510] = 18'b1010000101110111_10;
      patterns[511] = 18'b1011000101110111_11;
      patterns[512] = 18'b1000001000000000_00;
      patterns[513] = 18'b1001001000000000_01;
      patterns[514] = 18'b1010001000000000_10;
      patterns[515] = 18'b1011001000000000_11;
      patterns[516] = 18'b1000001000000001_00;
      patterns[517] = 18'b1001001000000001_01;
      patterns[518] = 18'b1010001000000001_10;
      patterns[519] = 18'b1011001000000001_11;
      patterns[520] = 18'b1000001000000010_00;
      patterns[521] = 18'b1001001000000010_01;
      patterns[522] = 18'b1010001000000010_10;
      patterns[523] = 18'b1011001000000010_11;
      patterns[524] = 18'b1000001000000011_00;
      patterns[525] = 18'b1001001000000011_01;
      patterns[526] = 18'b1010001000000011_10;
      patterns[527] = 18'b1011001000000011_11;
      patterns[528] = 18'b1000001000000100_00;
      patterns[529] = 18'b1001001000000100_01;
      patterns[530] = 18'b1010001000000100_10;
      patterns[531] = 18'b1011001000000100_11;
      patterns[532] = 18'b1000001000000101_00;
      patterns[533] = 18'b1001001000000101_01;
      patterns[534] = 18'b1010001000000101_10;
      patterns[535] = 18'b1011001000000101_11;
      patterns[536] = 18'b1000001000000110_00;
      patterns[537] = 18'b1001001000000110_01;
      patterns[538] = 18'b1010001000000110_10;
      patterns[539] = 18'b1011001000000110_11;
      patterns[540] = 18'b1000001000000111_00;
      patterns[541] = 18'b1001001000000111_01;
      patterns[542] = 18'b1010001000000111_10;
      patterns[543] = 18'b1011001000000111_11;
      patterns[544] = 18'b1000001000010000_00;
      patterns[545] = 18'b1001001000010000_01;
      patterns[546] = 18'b1010001000010000_10;
      patterns[547] = 18'b1011001000010000_11;
      patterns[548] = 18'b1000001000010001_00;
      patterns[549] = 18'b1001001000010001_01;
      patterns[550] = 18'b1010001000010001_10;
      patterns[551] = 18'b1011001000010001_11;
      patterns[552] = 18'b1000001000010010_00;
      patterns[553] = 18'b1001001000010010_01;
      patterns[554] = 18'b1010001000010010_10;
      patterns[555] = 18'b1011001000010010_11;
      patterns[556] = 18'b1000001000010011_00;
      patterns[557] = 18'b1001001000010011_01;
      patterns[558] = 18'b1010001000010011_10;
      patterns[559] = 18'b1011001000010011_11;
      patterns[560] = 18'b1000001000010100_00;
      patterns[561] = 18'b1001001000010100_01;
      patterns[562] = 18'b1010001000010100_10;
      patterns[563] = 18'b1011001000010100_11;
      patterns[564] = 18'b1000001000010101_00;
      patterns[565] = 18'b1001001000010101_01;
      patterns[566] = 18'b1010001000010101_10;
      patterns[567] = 18'b1011001000010101_11;
      patterns[568] = 18'b1000001000010110_00;
      patterns[569] = 18'b1001001000010110_01;
      patterns[570] = 18'b1010001000010110_10;
      patterns[571] = 18'b1011001000010110_11;
      patterns[572] = 18'b1000001000010111_00;
      patterns[573] = 18'b1001001000010111_01;
      patterns[574] = 18'b1010001000010111_10;
      patterns[575] = 18'b1011001000010111_11;
      patterns[576] = 18'b1000001000100000_00;
      patterns[577] = 18'b1001001000100000_01;
      patterns[578] = 18'b1010001000100000_10;
      patterns[579] = 18'b1011001000100000_11;
      patterns[580] = 18'b1000001000100001_00;
      patterns[581] = 18'b1001001000100001_01;
      patterns[582] = 18'b1010001000100001_10;
      patterns[583] = 18'b1011001000100001_11;
      patterns[584] = 18'b1000001000100010_00;
      patterns[585] = 18'b1001001000100010_01;
      patterns[586] = 18'b1010001000100010_10;
      patterns[587] = 18'b1011001000100010_11;
      patterns[588] = 18'b1000001000100011_00;
      patterns[589] = 18'b1001001000100011_01;
      patterns[590] = 18'b1010001000100011_10;
      patterns[591] = 18'b1011001000100011_11;
      patterns[592] = 18'b1000001000100100_00;
      patterns[593] = 18'b1001001000100100_01;
      patterns[594] = 18'b1010001000100100_10;
      patterns[595] = 18'b1011001000100100_11;
      patterns[596] = 18'b1000001000100101_00;
      patterns[597] = 18'b1001001000100101_01;
      patterns[598] = 18'b1010001000100101_10;
      patterns[599] = 18'b1011001000100101_11;
      patterns[600] = 18'b1000001000100110_00;
      patterns[601] = 18'b1001001000100110_01;
      patterns[602] = 18'b1010001000100110_10;
      patterns[603] = 18'b1011001000100110_11;
      patterns[604] = 18'b1000001000100111_00;
      patterns[605] = 18'b1001001000100111_01;
      patterns[606] = 18'b1010001000100111_10;
      patterns[607] = 18'b1011001000100111_11;
      patterns[608] = 18'b1000001000110000_00;
      patterns[609] = 18'b1001001000110000_01;
      patterns[610] = 18'b1010001000110000_10;
      patterns[611] = 18'b1011001000110000_11;
      patterns[612] = 18'b1000001000110001_00;
      patterns[613] = 18'b1001001000110001_01;
      patterns[614] = 18'b1010001000110001_10;
      patterns[615] = 18'b1011001000110001_11;
      patterns[616] = 18'b1000001000110010_00;
      patterns[617] = 18'b1001001000110010_01;
      patterns[618] = 18'b1010001000110010_10;
      patterns[619] = 18'b1011001000110010_11;
      patterns[620] = 18'b1000001000110011_00;
      patterns[621] = 18'b1001001000110011_01;
      patterns[622] = 18'b1010001000110011_10;
      patterns[623] = 18'b1011001000110011_11;
      patterns[624] = 18'b1000001000110100_00;
      patterns[625] = 18'b1001001000110100_01;
      patterns[626] = 18'b1010001000110100_10;
      patterns[627] = 18'b1011001000110100_11;
      patterns[628] = 18'b1000001000110101_00;
      patterns[629] = 18'b1001001000110101_01;
      patterns[630] = 18'b1010001000110101_10;
      patterns[631] = 18'b1011001000110101_11;
      patterns[632] = 18'b1000001000110110_00;
      patterns[633] = 18'b1001001000110110_01;
      patterns[634] = 18'b1010001000110110_10;
      patterns[635] = 18'b1011001000110110_11;
      patterns[636] = 18'b1000001000110111_00;
      patterns[637] = 18'b1001001000110111_01;
      patterns[638] = 18'b1010001000110111_10;
      patterns[639] = 18'b1011001000110111_11;
      patterns[640] = 18'b1000001001000000_00;
      patterns[641] = 18'b1001001001000000_01;
      patterns[642] = 18'b1010001001000000_10;
      patterns[643] = 18'b1011001001000000_11;
      patterns[644] = 18'b1000001001000001_00;
      patterns[645] = 18'b1001001001000001_01;
      patterns[646] = 18'b1010001001000001_10;
      patterns[647] = 18'b1011001001000001_11;
      patterns[648] = 18'b1000001001000010_00;
      patterns[649] = 18'b1001001001000010_01;
      patterns[650] = 18'b1010001001000010_10;
      patterns[651] = 18'b1011001001000010_11;
      patterns[652] = 18'b1000001001000011_00;
      patterns[653] = 18'b1001001001000011_01;
      patterns[654] = 18'b1010001001000011_10;
      patterns[655] = 18'b1011001001000011_11;
      patterns[656] = 18'b1000001001000100_00;
      patterns[657] = 18'b1001001001000100_01;
      patterns[658] = 18'b1010001001000100_10;
      patterns[659] = 18'b1011001001000100_11;
      patterns[660] = 18'b1000001001000101_00;
      patterns[661] = 18'b1001001001000101_01;
      patterns[662] = 18'b1010001001000101_10;
      patterns[663] = 18'b1011001001000101_11;
      patterns[664] = 18'b1000001001000110_00;
      patterns[665] = 18'b1001001001000110_01;
      patterns[666] = 18'b1010001001000110_10;
      patterns[667] = 18'b1011001001000110_11;
      patterns[668] = 18'b1000001001000111_00;
      patterns[669] = 18'b1001001001000111_01;
      patterns[670] = 18'b1010001001000111_10;
      patterns[671] = 18'b1011001001000111_11;
      patterns[672] = 18'b1000001001010000_00;
      patterns[673] = 18'b1001001001010000_01;
      patterns[674] = 18'b1010001001010000_10;
      patterns[675] = 18'b1011001001010000_11;
      patterns[676] = 18'b1000001001010001_00;
      patterns[677] = 18'b1001001001010001_01;
      patterns[678] = 18'b1010001001010001_10;
      patterns[679] = 18'b1011001001010001_11;
      patterns[680] = 18'b1000001001010010_00;
      patterns[681] = 18'b1001001001010010_01;
      patterns[682] = 18'b1010001001010010_10;
      patterns[683] = 18'b1011001001010010_11;
      patterns[684] = 18'b1000001001010011_00;
      patterns[685] = 18'b1001001001010011_01;
      patterns[686] = 18'b1010001001010011_10;
      patterns[687] = 18'b1011001001010011_11;
      patterns[688] = 18'b1000001001010100_00;
      patterns[689] = 18'b1001001001010100_01;
      patterns[690] = 18'b1010001001010100_10;
      patterns[691] = 18'b1011001001010100_11;
      patterns[692] = 18'b1000001001010101_00;
      patterns[693] = 18'b1001001001010101_01;
      patterns[694] = 18'b1010001001010101_10;
      patterns[695] = 18'b1011001001010101_11;
      patterns[696] = 18'b1000001001010110_00;
      patterns[697] = 18'b1001001001010110_01;
      patterns[698] = 18'b1010001001010110_10;
      patterns[699] = 18'b1011001001010110_11;
      patterns[700] = 18'b1000001001010111_00;
      patterns[701] = 18'b1001001001010111_01;
      patterns[702] = 18'b1010001001010111_10;
      patterns[703] = 18'b1011001001010111_11;
      patterns[704] = 18'b1000001001100000_00;
      patterns[705] = 18'b1001001001100000_01;
      patterns[706] = 18'b1010001001100000_10;
      patterns[707] = 18'b1011001001100000_11;
      patterns[708] = 18'b1000001001100001_00;
      patterns[709] = 18'b1001001001100001_01;
      patterns[710] = 18'b1010001001100001_10;
      patterns[711] = 18'b1011001001100001_11;
      patterns[712] = 18'b1000001001100010_00;
      patterns[713] = 18'b1001001001100010_01;
      patterns[714] = 18'b1010001001100010_10;
      patterns[715] = 18'b1011001001100010_11;
      patterns[716] = 18'b1000001001100011_00;
      patterns[717] = 18'b1001001001100011_01;
      patterns[718] = 18'b1010001001100011_10;
      patterns[719] = 18'b1011001001100011_11;
      patterns[720] = 18'b1000001001100100_00;
      patterns[721] = 18'b1001001001100100_01;
      patterns[722] = 18'b1010001001100100_10;
      patterns[723] = 18'b1011001001100100_11;
      patterns[724] = 18'b1000001001100101_00;
      patterns[725] = 18'b1001001001100101_01;
      patterns[726] = 18'b1010001001100101_10;
      patterns[727] = 18'b1011001001100101_11;
      patterns[728] = 18'b1000001001100110_00;
      patterns[729] = 18'b1001001001100110_01;
      patterns[730] = 18'b1010001001100110_10;
      patterns[731] = 18'b1011001001100110_11;
      patterns[732] = 18'b1000001001100111_00;
      patterns[733] = 18'b1001001001100111_01;
      patterns[734] = 18'b1010001001100111_10;
      patterns[735] = 18'b1011001001100111_11;
      patterns[736] = 18'b1000001001110000_00;
      patterns[737] = 18'b1001001001110000_01;
      patterns[738] = 18'b1010001001110000_10;
      patterns[739] = 18'b1011001001110000_11;
      patterns[740] = 18'b1000001001110001_00;
      patterns[741] = 18'b1001001001110001_01;
      patterns[742] = 18'b1010001001110001_10;
      patterns[743] = 18'b1011001001110001_11;
      patterns[744] = 18'b1000001001110010_00;
      patterns[745] = 18'b1001001001110010_01;
      patterns[746] = 18'b1010001001110010_10;
      patterns[747] = 18'b1011001001110010_11;
      patterns[748] = 18'b1000001001110011_00;
      patterns[749] = 18'b1001001001110011_01;
      patterns[750] = 18'b1010001001110011_10;
      patterns[751] = 18'b1011001001110011_11;
      patterns[752] = 18'b1000001001110100_00;
      patterns[753] = 18'b1001001001110100_01;
      patterns[754] = 18'b1010001001110100_10;
      patterns[755] = 18'b1011001001110100_11;
      patterns[756] = 18'b1000001001110101_00;
      patterns[757] = 18'b1001001001110101_01;
      patterns[758] = 18'b1010001001110101_10;
      patterns[759] = 18'b1011001001110101_11;
      patterns[760] = 18'b1000001001110110_00;
      patterns[761] = 18'b1001001001110110_01;
      patterns[762] = 18'b1010001001110110_10;
      patterns[763] = 18'b1011001001110110_11;
      patterns[764] = 18'b1000001001110111_00;
      patterns[765] = 18'b1001001001110111_01;
      patterns[766] = 18'b1010001001110111_10;
      patterns[767] = 18'b1011001001110111_11;
      patterns[768] = 18'b1000001100000000_00;
      patterns[769] = 18'b1001001100000000_01;
      patterns[770] = 18'b1010001100000000_10;
      patterns[771] = 18'b1011001100000000_11;
      patterns[772] = 18'b1000001100000001_00;
      patterns[773] = 18'b1001001100000001_01;
      patterns[774] = 18'b1010001100000001_10;
      patterns[775] = 18'b1011001100000001_11;
      patterns[776] = 18'b1000001100000010_00;
      patterns[777] = 18'b1001001100000010_01;
      patterns[778] = 18'b1010001100000010_10;
      patterns[779] = 18'b1011001100000010_11;
      patterns[780] = 18'b1000001100000011_00;
      patterns[781] = 18'b1001001100000011_01;
      patterns[782] = 18'b1010001100000011_10;
      patterns[783] = 18'b1011001100000011_11;
      patterns[784] = 18'b1000001100000100_00;
      patterns[785] = 18'b1001001100000100_01;
      patterns[786] = 18'b1010001100000100_10;
      patterns[787] = 18'b1011001100000100_11;
      patterns[788] = 18'b1000001100000101_00;
      patterns[789] = 18'b1001001100000101_01;
      patterns[790] = 18'b1010001100000101_10;
      patterns[791] = 18'b1011001100000101_11;
      patterns[792] = 18'b1000001100000110_00;
      patterns[793] = 18'b1001001100000110_01;
      patterns[794] = 18'b1010001100000110_10;
      patterns[795] = 18'b1011001100000110_11;
      patterns[796] = 18'b1000001100000111_00;
      patterns[797] = 18'b1001001100000111_01;
      patterns[798] = 18'b1010001100000111_10;
      patterns[799] = 18'b1011001100000111_11;
      patterns[800] = 18'b1000001100010000_00;
      patterns[801] = 18'b1001001100010000_01;
      patterns[802] = 18'b1010001100010000_10;
      patterns[803] = 18'b1011001100010000_11;
      patterns[804] = 18'b1000001100010001_00;
      patterns[805] = 18'b1001001100010001_01;
      patterns[806] = 18'b1010001100010001_10;
      patterns[807] = 18'b1011001100010001_11;
      patterns[808] = 18'b1000001100010010_00;
      patterns[809] = 18'b1001001100010010_01;
      patterns[810] = 18'b1010001100010010_10;
      patterns[811] = 18'b1011001100010010_11;
      patterns[812] = 18'b1000001100010011_00;
      patterns[813] = 18'b1001001100010011_01;
      patterns[814] = 18'b1010001100010011_10;
      patterns[815] = 18'b1011001100010011_11;
      patterns[816] = 18'b1000001100010100_00;
      patterns[817] = 18'b1001001100010100_01;
      patterns[818] = 18'b1010001100010100_10;
      patterns[819] = 18'b1011001100010100_11;
      patterns[820] = 18'b1000001100010101_00;
      patterns[821] = 18'b1001001100010101_01;
      patterns[822] = 18'b1010001100010101_10;
      patterns[823] = 18'b1011001100010101_11;
      patterns[824] = 18'b1000001100010110_00;
      patterns[825] = 18'b1001001100010110_01;
      patterns[826] = 18'b1010001100010110_10;
      patterns[827] = 18'b1011001100010110_11;
      patterns[828] = 18'b1000001100010111_00;
      patterns[829] = 18'b1001001100010111_01;
      patterns[830] = 18'b1010001100010111_10;
      patterns[831] = 18'b1011001100010111_11;
      patterns[832] = 18'b1000001100100000_00;
      patterns[833] = 18'b1001001100100000_01;
      patterns[834] = 18'b1010001100100000_10;
      patterns[835] = 18'b1011001100100000_11;
      patterns[836] = 18'b1000001100100001_00;
      patterns[837] = 18'b1001001100100001_01;
      patterns[838] = 18'b1010001100100001_10;
      patterns[839] = 18'b1011001100100001_11;
      patterns[840] = 18'b1000001100100010_00;
      patterns[841] = 18'b1001001100100010_01;
      patterns[842] = 18'b1010001100100010_10;
      patterns[843] = 18'b1011001100100010_11;
      patterns[844] = 18'b1000001100100011_00;
      patterns[845] = 18'b1001001100100011_01;
      patterns[846] = 18'b1010001100100011_10;
      patterns[847] = 18'b1011001100100011_11;
      patterns[848] = 18'b1000001100100100_00;
      patterns[849] = 18'b1001001100100100_01;
      patterns[850] = 18'b1010001100100100_10;
      patterns[851] = 18'b1011001100100100_11;
      patterns[852] = 18'b1000001100100101_00;
      patterns[853] = 18'b1001001100100101_01;
      patterns[854] = 18'b1010001100100101_10;
      patterns[855] = 18'b1011001100100101_11;
      patterns[856] = 18'b1000001100100110_00;
      patterns[857] = 18'b1001001100100110_01;
      patterns[858] = 18'b1010001100100110_10;
      patterns[859] = 18'b1011001100100110_11;
      patterns[860] = 18'b1000001100100111_00;
      patterns[861] = 18'b1001001100100111_01;
      patterns[862] = 18'b1010001100100111_10;
      patterns[863] = 18'b1011001100100111_11;
      patterns[864] = 18'b1000001100110000_00;
      patterns[865] = 18'b1001001100110000_01;
      patterns[866] = 18'b1010001100110000_10;
      patterns[867] = 18'b1011001100110000_11;
      patterns[868] = 18'b1000001100110001_00;
      patterns[869] = 18'b1001001100110001_01;
      patterns[870] = 18'b1010001100110001_10;
      patterns[871] = 18'b1011001100110001_11;
      patterns[872] = 18'b1000001100110010_00;
      patterns[873] = 18'b1001001100110010_01;
      patterns[874] = 18'b1010001100110010_10;
      patterns[875] = 18'b1011001100110010_11;
      patterns[876] = 18'b1000001100110011_00;
      patterns[877] = 18'b1001001100110011_01;
      patterns[878] = 18'b1010001100110011_10;
      patterns[879] = 18'b1011001100110011_11;
      patterns[880] = 18'b1000001100110100_00;
      patterns[881] = 18'b1001001100110100_01;
      patterns[882] = 18'b1010001100110100_10;
      patterns[883] = 18'b1011001100110100_11;
      patterns[884] = 18'b1000001100110101_00;
      patterns[885] = 18'b1001001100110101_01;
      patterns[886] = 18'b1010001100110101_10;
      patterns[887] = 18'b1011001100110101_11;
      patterns[888] = 18'b1000001100110110_00;
      patterns[889] = 18'b1001001100110110_01;
      patterns[890] = 18'b1010001100110110_10;
      patterns[891] = 18'b1011001100110110_11;
      patterns[892] = 18'b1000001100110111_00;
      patterns[893] = 18'b1001001100110111_01;
      patterns[894] = 18'b1010001100110111_10;
      patterns[895] = 18'b1011001100110111_11;
      patterns[896] = 18'b1000001101000000_00;
      patterns[897] = 18'b1001001101000000_01;
      patterns[898] = 18'b1010001101000000_10;
      patterns[899] = 18'b1011001101000000_11;
      patterns[900] = 18'b1000001101000001_00;
      patterns[901] = 18'b1001001101000001_01;
      patterns[902] = 18'b1010001101000001_10;
      patterns[903] = 18'b1011001101000001_11;
      patterns[904] = 18'b1000001101000010_00;
      patterns[905] = 18'b1001001101000010_01;
      patterns[906] = 18'b1010001101000010_10;
      patterns[907] = 18'b1011001101000010_11;
      patterns[908] = 18'b1000001101000011_00;
      patterns[909] = 18'b1001001101000011_01;
      patterns[910] = 18'b1010001101000011_10;
      patterns[911] = 18'b1011001101000011_11;
      patterns[912] = 18'b1000001101000100_00;
      patterns[913] = 18'b1001001101000100_01;
      patterns[914] = 18'b1010001101000100_10;
      patterns[915] = 18'b1011001101000100_11;
      patterns[916] = 18'b1000001101000101_00;
      patterns[917] = 18'b1001001101000101_01;
      patterns[918] = 18'b1010001101000101_10;
      patterns[919] = 18'b1011001101000101_11;
      patterns[920] = 18'b1000001101000110_00;
      patterns[921] = 18'b1001001101000110_01;
      patterns[922] = 18'b1010001101000110_10;
      patterns[923] = 18'b1011001101000110_11;
      patterns[924] = 18'b1000001101000111_00;
      patterns[925] = 18'b1001001101000111_01;
      patterns[926] = 18'b1010001101000111_10;
      patterns[927] = 18'b1011001101000111_11;
      patterns[928] = 18'b1000001101010000_00;
      patterns[929] = 18'b1001001101010000_01;
      patterns[930] = 18'b1010001101010000_10;
      patterns[931] = 18'b1011001101010000_11;
      patterns[932] = 18'b1000001101010001_00;
      patterns[933] = 18'b1001001101010001_01;
      patterns[934] = 18'b1010001101010001_10;
      patterns[935] = 18'b1011001101010001_11;
      patterns[936] = 18'b1000001101010010_00;
      patterns[937] = 18'b1001001101010010_01;
      patterns[938] = 18'b1010001101010010_10;
      patterns[939] = 18'b1011001101010010_11;
      patterns[940] = 18'b1000001101010011_00;
      patterns[941] = 18'b1001001101010011_01;
      patterns[942] = 18'b1010001101010011_10;
      patterns[943] = 18'b1011001101010011_11;
      patterns[944] = 18'b1000001101010100_00;
      patterns[945] = 18'b1001001101010100_01;
      patterns[946] = 18'b1010001101010100_10;
      patterns[947] = 18'b1011001101010100_11;
      patterns[948] = 18'b1000001101010101_00;
      patterns[949] = 18'b1001001101010101_01;
      patterns[950] = 18'b1010001101010101_10;
      patterns[951] = 18'b1011001101010101_11;
      patterns[952] = 18'b1000001101010110_00;
      patterns[953] = 18'b1001001101010110_01;
      patterns[954] = 18'b1010001101010110_10;
      patterns[955] = 18'b1011001101010110_11;
      patterns[956] = 18'b1000001101010111_00;
      patterns[957] = 18'b1001001101010111_01;
      patterns[958] = 18'b1010001101010111_10;
      patterns[959] = 18'b1011001101010111_11;
      patterns[960] = 18'b1000001101100000_00;
      patterns[961] = 18'b1001001101100000_01;
      patterns[962] = 18'b1010001101100000_10;
      patterns[963] = 18'b1011001101100000_11;
      patterns[964] = 18'b1000001101100001_00;
      patterns[965] = 18'b1001001101100001_01;
      patterns[966] = 18'b1010001101100001_10;
      patterns[967] = 18'b1011001101100001_11;
      patterns[968] = 18'b1000001101100010_00;
      patterns[969] = 18'b1001001101100010_01;
      patterns[970] = 18'b1010001101100010_10;
      patterns[971] = 18'b1011001101100010_11;
      patterns[972] = 18'b1000001101100011_00;
      patterns[973] = 18'b1001001101100011_01;
      patterns[974] = 18'b1010001101100011_10;
      patterns[975] = 18'b1011001101100011_11;
      patterns[976] = 18'b1000001101100100_00;
      patterns[977] = 18'b1001001101100100_01;
      patterns[978] = 18'b1010001101100100_10;
      patterns[979] = 18'b1011001101100100_11;
      patterns[980] = 18'b1000001101100101_00;
      patterns[981] = 18'b1001001101100101_01;
      patterns[982] = 18'b1010001101100101_10;
      patterns[983] = 18'b1011001101100101_11;
      patterns[984] = 18'b1000001101100110_00;
      patterns[985] = 18'b1001001101100110_01;
      patterns[986] = 18'b1010001101100110_10;
      patterns[987] = 18'b1011001101100110_11;
      patterns[988] = 18'b1000001101100111_00;
      patterns[989] = 18'b1001001101100111_01;
      patterns[990] = 18'b1010001101100111_10;
      patterns[991] = 18'b1011001101100111_11;
      patterns[992] = 18'b1000001101110000_00;
      patterns[993] = 18'b1001001101110000_01;
      patterns[994] = 18'b1010001101110000_10;
      patterns[995] = 18'b1011001101110000_11;
      patterns[996] = 18'b1000001101110001_00;
      patterns[997] = 18'b1001001101110001_01;
      patterns[998] = 18'b1010001101110001_10;
      patterns[999] = 18'b1011001101110001_11;
      patterns[1000] = 18'b1000001101110010_00;
      patterns[1001] = 18'b1001001101110010_01;
      patterns[1002] = 18'b1010001101110010_10;
      patterns[1003] = 18'b1011001101110010_11;
      patterns[1004] = 18'b1000001101110011_00;
      patterns[1005] = 18'b1001001101110011_01;
      patterns[1006] = 18'b1010001101110011_10;
      patterns[1007] = 18'b1011001101110011_11;
      patterns[1008] = 18'b1000001101110100_00;
      patterns[1009] = 18'b1001001101110100_01;
      patterns[1010] = 18'b1010001101110100_10;
      patterns[1011] = 18'b1011001101110100_11;
      patterns[1012] = 18'b1000001101110101_00;
      patterns[1013] = 18'b1001001101110101_01;
      patterns[1014] = 18'b1010001101110101_10;
      patterns[1015] = 18'b1011001101110101_11;
      patterns[1016] = 18'b1000001101110110_00;
      patterns[1017] = 18'b1001001101110110_01;
      patterns[1018] = 18'b1010001101110110_10;
      patterns[1019] = 18'b1011001101110110_11;
      patterns[1020] = 18'b1000001101110111_00;
      patterns[1021] = 18'b1001001101110111_01;
      patterns[1022] = 18'b1010001101110111_10;
      patterns[1023] = 18'b1011001101110111_11;
      patterns[1024] = 18'b1000010000000000_00;
      patterns[1025] = 18'b1001010000000000_01;
      patterns[1026] = 18'b1010010000000000_10;
      patterns[1027] = 18'b1011010000000000_11;
      patterns[1028] = 18'b1000010000000001_00;
      patterns[1029] = 18'b1001010000000001_01;
      patterns[1030] = 18'b1010010000000001_10;
      patterns[1031] = 18'b1011010000000001_11;
      patterns[1032] = 18'b1000010000000010_00;
      patterns[1033] = 18'b1001010000000010_01;
      patterns[1034] = 18'b1010010000000010_10;
      patterns[1035] = 18'b1011010000000010_11;
      patterns[1036] = 18'b1000010000000011_00;
      patterns[1037] = 18'b1001010000000011_01;
      patterns[1038] = 18'b1010010000000011_10;
      patterns[1039] = 18'b1011010000000011_11;
      patterns[1040] = 18'b1000010000000100_00;
      patterns[1041] = 18'b1001010000000100_01;
      patterns[1042] = 18'b1010010000000100_10;
      patterns[1043] = 18'b1011010000000100_11;
      patterns[1044] = 18'b1000010000000101_00;
      patterns[1045] = 18'b1001010000000101_01;
      patterns[1046] = 18'b1010010000000101_10;
      patterns[1047] = 18'b1011010000000101_11;
      patterns[1048] = 18'b1000010000000110_00;
      patterns[1049] = 18'b1001010000000110_01;
      patterns[1050] = 18'b1010010000000110_10;
      patterns[1051] = 18'b1011010000000110_11;
      patterns[1052] = 18'b1000010000000111_00;
      patterns[1053] = 18'b1001010000000111_01;
      patterns[1054] = 18'b1010010000000111_10;
      patterns[1055] = 18'b1011010000000111_11;
      patterns[1056] = 18'b1000010000010000_00;
      patterns[1057] = 18'b1001010000010000_01;
      patterns[1058] = 18'b1010010000010000_10;
      patterns[1059] = 18'b1011010000010000_11;
      patterns[1060] = 18'b1000010000010001_00;
      patterns[1061] = 18'b1001010000010001_01;
      patterns[1062] = 18'b1010010000010001_10;
      patterns[1063] = 18'b1011010000010001_11;
      patterns[1064] = 18'b1000010000010010_00;
      patterns[1065] = 18'b1001010000010010_01;
      patterns[1066] = 18'b1010010000010010_10;
      patterns[1067] = 18'b1011010000010010_11;
      patterns[1068] = 18'b1000010000010011_00;
      patterns[1069] = 18'b1001010000010011_01;
      patterns[1070] = 18'b1010010000010011_10;
      patterns[1071] = 18'b1011010000010011_11;
      patterns[1072] = 18'b1000010000010100_00;
      patterns[1073] = 18'b1001010000010100_01;
      patterns[1074] = 18'b1010010000010100_10;
      patterns[1075] = 18'b1011010000010100_11;
      patterns[1076] = 18'b1000010000010101_00;
      patterns[1077] = 18'b1001010000010101_01;
      patterns[1078] = 18'b1010010000010101_10;
      patterns[1079] = 18'b1011010000010101_11;
      patterns[1080] = 18'b1000010000010110_00;
      patterns[1081] = 18'b1001010000010110_01;
      patterns[1082] = 18'b1010010000010110_10;
      patterns[1083] = 18'b1011010000010110_11;
      patterns[1084] = 18'b1000010000010111_00;
      patterns[1085] = 18'b1001010000010111_01;
      patterns[1086] = 18'b1010010000010111_10;
      patterns[1087] = 18'b1011010000010111_11;
      patterns[1088] = 18'b1000010000100000_00;
      patterns[1089] = 18'b1001010000100000_01;
      patterns[1090] = 18'b1010010000100000_10;
      patterns[1091] = 18'b1011010000100000_11;
      patterns[1092] = 18'b1000010000100001_00;
      patterns[1093] = 18'b1001010000100001_01;
      patterns[1094] = 18'b1010010000100001_10;
      patterns[1095] = 18'b1011010000100001_11;
      patterns[1096] = 18'b1000010000100010_00;
      patterns[1097] = 18'b1001010000100010_01;
      patterns[1098] = 18'b1010010000100010_10;
      patterns[1099] = 18'b1011010000100010_11;
      patterns[1100] = 18'b1000010000100011_00;
      patterns[1101] = 18'b1001010000100011_01;
      patterns[1102] = 18'b1010010000100011_10;
      patterns[1103] = 18'b1011010000100011_11;
      patterns[1104] = 18'b1000010000100100_00;
      patterns[1105] = 18'b1001010000100100_01;
      patterns[1106] = 18'b1010010000100100_10;
      patterns[1107] = 18'b1011010000100100_11;
      patterns[1108] = 18'b1000010000100101_00;
      patterns[1109] = 18'b1001010000100101_01;
      patterns[1110] = 18'b1010010000100101_10;
      patterns[1111] = 18'b1011010000100101_11;
      patterns[1112] = 18'b1000010000100110_00;
      patterns[1113] = 18'b1001010000100110_01;
      patterns[1114] = 18'b1010010000100110_10;
      patterns[1115] = 18'b1011010000100110_11;
      patterns[1116] = 18'b1000010000100111_00;
      patterns[1117] = 18'b1001010000100111_01;
      patterns[1118] = 18'b1010010000100111_10;
      patterns[1119] = 18'b1011010000100111_11;
      patterns[1120] = 18'b1000010000110000_00;
      patterns[1121] = 18'b1001010000110000_01;
      patterns[1122] = 18'b1010010000110000_10;
      patterns[1123] = 18'b1011010000110000_11;
      patterns[1124] = 18'b1000010000110001_00;
      patterns[1125] = 18'b1001010000110001_01;
      patterns[1126] = 18'b1010010000110001_10;
      patterns[1127] = 18'b1011010000110001_11;
      patterns[1128] = 18'b1000010000110010_00;
      patterns[1129] = 18'b1001010000110010_01;
      patterns[1130] = 18'b1010010000110010_10;
      patterns[1131] = 18'b1011010000110010_11;
      patterns[1132] = 18'b1000010000110011_00;
      patterns[1133] = 18'b1001010000110011_01;
      patterns[1134] = 18'b1010010000110011_10;
      patterns[1135] = 18'b1011010000110011_11;
      patterns[1136] = 18'b1000010000110100_00;
      patterns[1137] = 18'b1001010000110100_01;
      patterns[1138] = 18'b1010010000110100_10;
      patterns[1139] = 18'b1011010000110100_11;
      patterns[1140] = 18'b1000010000110101_00;
      patterns[1141] = 18'b1001010000110101_01;
      patterns[1142] = 18'b1010010000110101_10;
      patterns[1143] = 18'b1011010000110101_11;
      patterns[1144] = 18'b1000010000110110_00;
      patterns[1145] = 18'b1001010000110110_01;
      patterns[1146] = 18'b1010010000110110_10;
      patterns[1147] = 18'b1011010000110110_11;
      patterns[1148] = 18'b1000010000110111_00;
      patterns[1149] = 18'b1001010000110111_01;
      patterns[1150] = 18'b1010010000110111_10;
      patterns[1151] = 18'b1011010000110111_11;
      patterns[1152] = 18'b1000010001000000_00;
      patterns[1153] = 18'b1001010001000000_01;
      patterns[1154] = 18'b1010010001000000_10;
      patterns[1155] = 18'b1011010001000000_11;
      patterns[1156] = 18'b1000010001000001_00;
      patterns[1157] = 18'b1001010001000001_01;
      patterns[1158] = 18'b1010010001000001_10;
      patterns[1159] = 18'b1011010001000001_11;
      patterns[1160] = 18'b1000010001000010_00;
      patterns[1161] = 18'b1001010001000010_01;
      patterns[1162] = 18'b1010010001000010_10;
      patterns[1163] = 18'b1011010001000010_11;
      patterns[1164] = 18'b1000010001000011_00;
      patterns[1165] = 18'b1001010001000011_01;
      patterns[1166] = 18'b1010010001000011_10;
      patterns[1167] = 18'b1011010001000011_11;
      patterns[1168] = 18'b1000010001000100_00;
      patterns[1169] = 18'b1001010001000100_01;
      patterns[1170] = 18'b1010010001000100_10;
      patterns[1171] = 18'b1011010001000100_11;
      patterns[1172] = 18'b1000010001000101_00;
      patterns[1173] = 18'b1001010001000101_01;
      patterns[1174] = 18'b1010010001000101_10;
      patterns[1175] = 18'b1011010001000101_11;
      patterns[1176] = 18'b1000010001000110_00;
      patterns[1177] = 18'b1001010001000110_01;
      patterns[1178] = 18'b1010010001000110_10;
      patterns[1179] = 18'b1011010001000110_11;
      patterns[1180] = 18'b1000010001000111_00;
      patterns[1181] = 18'b1001010001000111_01;
      patterns[1182] = 18'b1010010001000111_10;
      patterns[1183] = 18'b1011010001000111_11;
      patterns[1184] = 18'b1000010001010000_00;
      patterns[1185] = 18'b1001010001010000_01;
      patterns[1186] = 18'b1010010001010000_10;
      patterns[1187] = 18'b1011010001010000_11;
      patterns[1188] = 18'b1000010001010001_00;
      patterns[1189] = 18'b1001010001010001_01;
      patterns[1190] = 18'b1010010001010001_10;
      patterns[1191] = 18'b1011010001010001_11;
      patterns[1192] = 18'b1000010001010010_00;
      patterns[1193] = 18'b1001010001010010_01;
      patterns[1194] = 18'b1010010001010010_10;
      patterns[1195] = 18'b1011010001010010_11;
      patterns[1196] = 18'b1000010001010011_00;
      patterns[1197] = 18'b1001010001010011_01;
      patterns[1198] = 18'b1010010001010011_10;
      patterns[1199] = 18'b1011010001010011_11;
      patterns[1200] = 18'b1000010001010100_00;
      patterns[1201] = 18'b1001010001010100_01;
      patterns[1202] = 18'b1010010001010100_10;
      patterns[1203] = 18'b1011010001010100_11;
      patterns[1204] = 18'b1000010001010101_00;
      patterns[1205] = 18'b1001010001010101_01;
      patterns[1206] = 18'b1010010001010101_10;
      patterns[1207] = 18'b1011010001010101_11;
      patterns[1208] = 18'b1000010001010110_00;
      patterns[1209] = 18'b1001010001010110_01;
      patterns[1210] = 18'b1010010001010110_10;
      patterns[1211] = 18'b1011010001010110_11;
      patterns[1212] = 18'b1000010001010111_00;
      patterns[1213] = 18'b1001010001010111_01;
      patterns[1214] = 18'b1010010001010111_10;
      patterns[1215] = 18'b1011010001010111_11;
      patterns[1216] = 18'b1000010001100000_00;
      patterns[1217] = 18'b1001010001100000_01;
      patterns[1218] = 18'b1010010001100000_10;
      patterns[1219] = 18'b1011010001100000_11;
      patterns[1220] = 18'b1000010001100001_00;
      patterns[1221] = 18'b1001010001100001_01;
      patterns[1222] = 18'b1010010001100001_10;
      patterns[1223] = 18'b1011010001100001_11;
      patterns[1224] = 18'b1000010001100010_00;
      patterns[1225] = 18'b1001010001100010_01;
      patterns[1226] = 18'b1010010001100010_10;
      patterns[1227] = 18'b1011010001100010_11;
      patterns[1228] = 18'b1000010001100011_00;
      patterns[1229] = 18'b1001010001100011_01;
      patterns[1230] = 18'b1010010001100011_10;
      patterns[1231] = 18'b1011010001100011_11;
      patterns[1232] = 18'b1000010001100100_00;
      patterns[1233] = 18'b1001010001100100_01;
      patterns[1234] = 18'b1010010001100100_10;
      patterns[1235] = 18'b1011010001100100_11;
      patterns[1236] = 18'b1000010001100101_00;
      patterns[1237] = 18'b1001010001100101_01;
      patterns[1238] = 18'b1010010001100101_10;
      patterns[1239] = 18'b1011010001100101_11;
      patterns[1240] = 18'b1000010001100110_00;
      patterns[1241] = 18'b1001010001100110_01;
      patterns[1242] = 18'b1010010001100110_10;
      patterns[1243] = 18'b1011010001100110_11;
      patterns[1244] = 18'b1000010001100111_00;
      patterns[1245] = 18'b1001010001100111_01;
      patterns[1246] = 18'b1010010001100111_10;
      patterns[1247] = 18'b1011010001100111_11;
      patterns[1248] = 18'b1000010001110000_00;
      patterns[1249] = 18'b1001010001110000_01;
      patterns[1250] = 18'b1010010001110000_10;
      patterns[1251] = 18'b1011010001110000_11;
      patterns[1252] = 18'b1000010001110001_00;
      patterns[1253] = 18'b1001010001110001_01;
      patterns[1254] = 18'b1010010001110001_10;
      patterns[1255] = 18'b1011010001110001_11;
      patterns[1256] = 18'b1000010001110010_00;
      patterns[1257] = 18'b1001010001110010_01;
      patterns[1258] = 18'b1010010001110010_10;
      patterns[1259] = 18'b1011010001110010_11;
      patterns[1260] = 18'b1000010001110011_00;
      patterns[1261] = 18'b1001010001110011_01;
      patterns[1262] = 18'b1010010001110011_10;
      patterns[1263] = 18'b1011010001110011_11;
      patterns[1264] = 18'b1000010001110100_00;
      patterns[1265] = 18'b1001010001110100_01;
      patterns[1266] = 18'b1010010001110100_10;
      patterns[1267] = 18'b1011010001110100_11;
      patterns[1268] = 18'b1000010001110101_00;
      patterns[1269] = 18'b1001010001110101_01;
      patterns[1270] = 18'b1010010001110101_10;
      patterns[1271] = 18'b1011010001110101_11;
      patterns[1272] = 18'b1000010001110110_00;
      patterns[1273] = 18'b1001010001110110_01;
      patterns[1274] = 18'b1010010001110110_10;
      patterns[1275] = 18'b1011010001110110_11;
      patterns[1276] = 18'b1000010001110111_00;
      patterns[1277] = 18'b1001010001110111_01;
      patterns[1278] = 18'b1010010001110111_10;
      patterns[1279] = 18'b1011010001110111_11;
      patterns[1280] = 18'b1000010100000000_00;
      patterns[1281] = 18'b1001010100000000_01;
      patterns[1282] = 18'b1010010100000000_10;
      patterns[1283] = 18'b1011010100000000_11;
      patterns[1284] = 18'b1000010100000001_00;
      patterns[1285] = 18'b1001010100000001_01;
      patterns[1286] = 18'b1010010100000001_10;
      patterns[1287] = 18'b1011010100000001_11;
      patterns[1288] = 18'b1000010100000010_00;
      patterns[1289] = 18'b1001010100000010_01;
      patterns[1290] = 18'b1010010100000010_10;
      patterns[1291] = 18'b1011010100000010_11;
      patterns[1292] = 18'b1000010100000011_00;
      patterns[1293] = 18'b1001010100000011_01;
      patterns[1294] = 18'b1010010100000011_10;
      patterns[1295] = 18'b1011010100000011_11;
      patterns[1296] = 18'b1000010100000100_00;
      patterns[1297] = 18'b1001010100000100_01;
      patterns[1298] = 18'b1010010100000100_10;
      patterns[1299] = 18'b1011010100000100_11;
      patterns[1300] = 18'b1000010100000101_00;
      patterns[1301] = 18'b1001010100000101_01;
      patterns[1302] = 18'b1010010100000101_10;
      patterns[1303] = 18'b1011010100000101_11;
      patterns[1304] = 18'b1000010100000110_00;
      patterns[1305] = 18'b1001010100000110_01;
      patterns[1306] = 18'b1010010100000110_10;
      patterns[1307] = 18'b1011010100000110_11;
      patterns[1308] = 18'b1000010100000111_00;
      patterns[1309] = 18'b1001010100000111_01;
      patterns[1310] = 18'b1010010100000111_10;
      patterns[1311] = 18'b1011010100000111_11;
      patterns[1312] = 18'b1000010100010000_00;
      patterns[1313] = 18'b1001010100010000_01;
      patterns[1314] = 18'b1010010100010000_10;
      patterns[1315] = 18'b1011010100010000_11;
      patterns[1316] = 18'b1000010100010001_00;
      patterns[1317] = 18'b1001010100010001_01;
      patterns[1318] = 18'b1010010100010001_10;
      patterns[1319] = 18'b1011010100010001_11;
      patterns[1320] = 18'b1000010100010010_00;
      patterns[1321] = 18'b1001010100010010_01;
      patterns[1322] = 18'b1010010100010010_10;
      patterns[1323] = 18'b1011010100010010_11;
      patterns[1324] = 18'b1000010100010011_00;
      patterns[1325] = 18'b1001010100010011_01;
      patterns[1326] = 18'b1010010100010011_10;
      patterns[1327] = 18'b1011010100010011_11;
      patterns[1328] = 18'b1000010100010100_00;
      patterns[1329] = 18'b1001010100010100_01;
      patterns[1330] = 18'b1010010100010100_10;
      patterns[1331] = 18'b1011010100010100_11;
      patterns[1332] = 18'b1000010100010101_00;
      patterns[1333] = 18'b1001010100010101_01;
      patterns[1334] = 18'b1010010100010101_10;
      patterns[1335] = 18'b1011010100010101_11;
      patterns[1336] = 18'b1000010100010110_00;
      patterns[1337] = 18'b1001010100010110_01;
      patterns[1338] = 18'b1010010100010110_10;
      patterns[1339] = 18'b1011010100010110_11;
      patterns[1340] = 18'b1000010100010111_00;
      patterns[1341] = 18'b1001010100010111_01;
      patterns[1342] = 18'b1010010100010111_10;
      patterns[1343] = 18'b1011010100010111_11;
      patterns[1344] = 18'b1000010100100000_00;
      patterns[1345] = 18'b1001010100100000_01;
      patterns[1346] = 18'b1010010100100000_10;
      patterns[1347] = 18'b1011010100100000_11;
      patterns[1348] = 18'b1000010100100001_00;
      patterns[1349] = 18'b1001010100100001_01;
      patterns[1350] = 18'b1010010100100001_10;
      patterns[1351] = 18'b1011010100100001_11;
      patterns[1352] = 18'b1000010100100010_00;
      patterns[1353] = 18'b1001010100100010_01;
      patterns[1354] = 18'b1010010100100010_10;
      patterns[1355] = 18'b1011010100100010_11;
      patterns[1356] = 18'b1000010100100011_00;
      patterns[1357] = 18'b1001010100100011_01;
      patterns[1358] = 18'b1010010100100011_10;
      patterns[1359] = 18'b1011010100100011_11;
      patterns[1360] = 18'b1000010100100100_00;
      patterns[1361] = 18'b1001010100100100_01;
      patterns[1362] = 18'b1010010100100100_10;
      patterns[1363] = 18'b1011010100100100_11;
      patterns[1364] = 18'b1000010100100101_00;
      patterns[1365] = 18'b1001010100100101_01;
      patterns[1366] = 18'b1010010100100101_10;
      patterns[1367] = 18'b1011010100100101_11;
      patterns[1368] = 18'b1000010100100110_00;
      patterns[1369] = 18'b1001010100100110_01;
      patterns[1370] = 18'b1010010100100110_10;
      patterns[1371] = 18'b1011010100100110_11;
      patterns[1372] = 18'b1000010100100111_00;
      patterns[1373] = 18'b1001010100100111_01;
      patterns[1374] = 18'b1010010100100111_10;
      patterns[1375] = 18'b1011010100100111_11;
      patterns[1376] = 18'b1000010100110000_00;
      patterns[1377] = 18'b1001010100110000_01;
      patterns[1378] = 18'b1010010100110000_10;
      patterns[1379] = 18'b1011010100110000_11;
      patterns[1380] = 18'b1000010100110001_00;
      patterns[1381] = 18'b1001010100110001_01;
      patterns[1382] = 18'b1010010100110001_10;
      patterns[1383] = 18'b1011010100110001_11;
      patterns[1384] = 18'b1000010100110010_00;
      patterns[1385] = 18'b1001010100110010_01;
      patterns[1386] = 18'b1010010100110010_10;
      patterns[1387] = 18'b1011010100110010_11;
      patterns[1388] = 18'b1000010100110011_00;
      patterns[1389] = 18'b1001010100110011_01;
      patterns[1390] = 18'b1010010100110011_10;
      patterns[1391] = 18'b1011010100110011_11;
      patterns[1392] = 18'b1000010100110100_00;
      patterns[1393] = 18'b1001010100110100_01;
      patterns[1394] = 18'b1010010100110100_10;
      patterns[1395] = 18'b1011010100110100_11;
      patterns[1396] = 18'b1000010100110101_00;
      patterns[1397] = 18'b1001010100110101_01;
      patterns[1398] = 18'b1010010100110101_10;
      patterns[1399] = 18'b1011010100110101_11;
      patterns[1400] = 18'b1000010100110110_00;
      patterns[1401] = 18'b1001010100110110_01;
      patterns[1402] = 18'b1010010100110110_10;
      patterns[1403] = 18'b1011010100110110_11;
      patterns[1404] = 18'b1000010100110111_00;
      patterns[1405] = 18'b1001010100110111_01;
      patterns[1406] = 18'b1010010100110111_10;
      patterns[1407] = 18'b1011010100110111_11;
      patterns[1408] = 18'b1000010101000000_00;
      patterns[1409] = 18'b1001010101000000_01;
      patterns[1410] = 18'b1010010101000000_10;
      patterns[1411] = 18'b1011010101000000_11;
      patterns[1412] = 18'b1000010101000001_00;
      patterns[1413] = 18'b1001010101000001_01;
      patterns[1414] = 18'b1010010101000001_10;
      patterns[1415] = 18'b1011010101000001_11;
      patterns[1416] = 18'b1000010101000010_00;
      patterns[1417] = 18'b1001010101000010_01;
      patterns[1418] = 18'b1010010101000010_10;
      patterns[1419] = 18'b1011010101000010_11;
      patterns[1420] = 18'b1000010101000011_00;
      patterns[1421] = 18'b1001010101000011_01;
      patterns[1422] = 18'b1010010101000011_10;
      patterns[1423] = 18'b1011010101000011_11;
      patterns[1424] = 18'b1000010101000100_00;
      patterns[1425] = 18'b1001010101000100_01;
      patterns[1426] = 18'b1010010101000100_10;
      patterns[1427] = 18'b1011010101000100_11;
      patterns[1428] = 18'b1000010101000101_00;
      patterns[1429] = 18'b1001010101000101_01;
      patterns[1430] = 18'b1010010101000101_10;
      patterns[1431] = 18'b1011010101000101_11;
      patterns[1432] = 18'b1000010101000110_00;
      patterns[1433] = 18'b1001010101000110_01;
      patterns[1434] = 18'b1010010101000110_10;
      patterns[1435] = 18'b1011010101000110_11;
      patterns[1436] = 18'b1000010101000111_00;
      patterns[1437] = 18'b1001010101000111_01;
      patterns[1438] = 18'b1010010101000111_10;
      patterns[1439] = 18'b1011010101000111_11;
      patterns[1440] = 18'b1000010101010000_00;
      patterns[1441] = 18'b1001010101010000_01;
      patterns[1442] = 18'b1010010101010000_10;
      patterns[1443] = 18'b1011010101010000_11;
      patterns[1444] = 18'b1000010101010001_00;
      patterns[1445] = 18'b1001010101010001_01;
      patterns[1446] = 18'b1010010101010001_10;
      patterns[1447] = 18'b1011010101010001_11;
      patterns[1448] = 18'b1000010101010010_00;
      patterns[1449] = 18'b1001010101010010_01;
      patterns[1450] = 18'b1010010101010010_10;
      patterns[1451] = 18'b1011010101010010_11;
      patterns[1452] = 18'b1000010101010011_00;
      patterns[1453] = 18'b1001010101010011_01;
      patterns[1454] = 18'b1010010101010011_10;
      patterns[1455] = 18'b1011010101010011_11;
      patterns[1456] = 18'b1000010101010100_00;
      patterns[1457] = 18'b1001010101010100_01;
      patterns[1458] = 18'b1010010101010100_10;
      patterns[1459] = 18'b1011010101010100_11;
      patterns[1460] = 18'b1000010101010101_00;
      patterns[1461] = 18'b1001010101010101_01;
      patterns[1462] = 18'b1010010101010101_10;
      patterns[1463] = 18'b1011010101010101_11;
      patterns[1464] = 18'b1000010101010110_00;
      patterns[1465] = 18'b1001010101010110_01;
      patterns[1466] = 18'b1010010101010110_10;
      patterns[1467] = 18'b1011010101010110_11;
      patterns[1468] = 18'b1000010101010111_00;
      patterns[1469] = 18'b1001010101010111_01;
      patterns[1470] = 18'b1010010101010111_10;
      patterns[1471] = 18'b1011010101010111_11;
      patterns[1472] = 18'b1000010101100000_00;
      patterns[1473] = 18'b1001010101100000_01;
      patterns[1474] = 18'b1010010101100000_10;
      patterns[1475] = 18'b1011010101100000_11;
      patterns[1476] = 18'b1000010101100001_00;
      patterns[1477] = 18'b1001010101100001_01;
      patterns[1478] = 18'b1010010101100001_10;
      patterns[1479] = 18'b1011010101100001_11;
      patterns[1480] = 18'b1000010101100010_00;
      patterns[1481] = 18'b1001010101100010_01;
      patterns[1482] = 18'b1010010101100010_10;
      patterns[1483] = 18'b1011010101100010_11;
      patterns[1484] = 18'b1000010101100011_00;
      patterns[1485] = 18'b1001010101100011_01;
      patterns[1486] = 18'b1010010101100011_10;
      patterns[1487] = 18'b1011010101100011_11;
      patterns[1488] = 18'b1000010101100100_00;
      patterns[1489] = 18'b1001010101100100_01;
      patterns[1490] = 18'b1010010101100100_10;
      patterns[1491] = 18'b1011010101100100_11;
      patterns[1492] = 18'b1000010101100101_00;
      patterns[1493] = 18'b1001010101100101_01;
      patterns[1494] = 18'b1010010101100101_10;
      patterns[1495] = 18'b1011010101100101_11;
      patterns[1496] = 18'b1000010101100110_00;
      patterns[1497] = 18'b1001010101100110_01;
      patterns[1498] = 18'b1010010101100110_10;
      patterns[1499] = 18'b1011010101100110_11;
      patterns[1500] = 18'b1000010101100111_00;
      patterns[1501] = 18'b1001010101100111_01;
      patterns[1502] = 18'b1010010101100111_10;
      patterns[1503] = 18'b1011010101100111_11;
      patterns[1504] = 18'b1000010101110000_00;
      patterns[1505] = 18'b1001010101110000_01;
      patterns[1506] = 18'b1010010101110000_10;
      patterns[1507] = 18'b1011010101110000_11;
      patterns[1508] = 18'b1000010101110001_00;
      patterns[1509] = 18'b1001010101110001_01;
      patterns[1510] = 18'b1010010101110001_10;
      patterns[1511] = 18'b1011010101110001_11;
      patterns[1512] = 18'b1000010101110010_00;
      patterns[1513] = 18'b1001010101110010_01;
      patterns[1514] = 18'b1010010101110010_10;
      patterns[1515] = 18'b1011010101110010_11;
      patterns[1516] = 18'b1000010101110011_00;
      patterns[1517] = 18'b1001010101110011_01;
      patterns[1518] = 18'b1010010101110011_10;
      patterns[1519] = 18'b1011010101110011_11;
      patterns[1520] = 18'b1000010101110100_00;
      patterns[1521] = 18'b1001010101110100_01;
      patterns[1522] = 18'b1010010101110100_10;
      patterns[1523] = 18'b1011010101110100_11;
      patterns[1524] = 18'b1000010101110101_00;
      patterns[1525] = 18'b1001010101110101_01;
      patterns[1526] = 18'b1010010101110101_10;
      patterns[1527] = 18'b1011010101110101_11;
      patterns[1528] = 18'b1000010101110110_00;
      patterns[1529] = 18'b1001010101110110_01;
      patterns[1530] = 18'b1010010101110110_10;
      patterns[1531] = 18'b1011010101110110_11;
      patterns[1532] = 18'b1000010101110111_00;
      patterns[1533] = 18'b1001010101110111_01;
      patterns[1534] = 18'b1010010101110111_10;
      patterns[1535] = 18'b1011010101110111_11;
      patterns[1536] = 18'b1000011000000000_00;
      patterns[1537] = 18'b1001011000000000_01;
      patterns[1538] = 18'b1010011000000000_10;
      patterns[1539] = 18'b1011011000000000_11;
      patterns[1540] = 18'b1000011000000001_00;
      patterns[1541] = 18'b1001011000000001_01;
      patterns[1542] = 18'b1010011000000001_10;
      patterns[1543] = 18'b1011011000000001_11;
      patterns[1544] = 18'b1000011000000010_00;
      patterns[1545] = 18'b1001011000000010_01;
      patterns[1546] = 18'b1010011000000010_10;
      patterns[1547] = 18'b1011011000000010_11;
      patterns[1548] = 18'b1000011000000011_00;
      patterns[1549] = 18'b1001011000000011_01;
      patterns[1550] = 18'b1010011000000011_10;
      patterns[1551] = 18'b1011011000000011_11;
      patterns[1552] = 18'b1000011000000100_00;
      patterns[1553] = 18'b1001011000000100_01;
      patterns[1554] = 18'b1010011000000100_10;
      patterns[1555] = 18'b1011011000000100_11;
      patterns[1556] = 18'b1000011000000101_00;
      patterns[1557] = 18'b1001011000000101_01;
      patterns[1558] = 18'b1010011000000101_10;
      patterns[1559] = 18'b1011011000000101_11;
      patterns[1560] = 18'b1000011000000110_00;
      patterns[1561] = 18'b1001011000000110_01;
      patterns[1562] = 18'b1010011000000110_10;
      patterns[1563] = 18'b1011011000000110_11;
      patterns[1564] = 18'b1000011000000111_00;
      patterns[1565] = 18'b1001011000000111_01;
      patterns[1566] = 18'b1010011000000111_10;
      patterns[1567] = 18'b1011011000000111_11;
      patterns[1568] = 18'b1000011000010000_00;
      patterns[1569] = 18'b1001011000010000_01;
      patterns[1570] = 18'b1010011000010000_10;
      patterns[1571] = 18'b1011011000010000_11;
      patterns[1572] = 18'b1000011000010001_00;
      patterns[1573] = 18'b1001011000010001_01;
      patterns[1574] = 18'b1010011000010001_10;
      patterns[1575] = 18'b1011011000010001_11;
      patterns[1576] = 18'b1000011000010010_00;
      patterns[1577] = 18'b1001011000010010_01;
      patterns[1578] = 18'b1010011000010010_10;
      patterns[1579] = 18'b1011011000010010_11;
      patterns[1580] = 18'b1000011000010011_00;
      patterns[1581] = 18'b1001011000010011_01;
      patterns[1582] = 18'b1010011000010011_10;
      patterns[1583] = 18'b1011011000010011_11;
      patterns[1584] = 18'b1000011000010100_00;
      patterns[1585] = 18'b1001011000010100_01;
      patterns[1586] = 18'b1010011000010100_10;
      patterns[1587] = 18'b1011011000010100_11;
      patterns[1588] = 18'b1000011000010101_00;
      patterns[1589] = 18'b1001011000010101_01;
      patterns[1590] = 18'b1010011000010101_10;
      patterns[1591] = 18'b1011011000010101_11;
      patterns[1592] = 18'b1000011000010110_00;
      patterns[1593] = 18'b1001011000010110_01;
      patterns[1594] = 18'b1010011000010110_10;
      patterns[1595] = 18'b1011011000010110_11;
      patterns[1596] = 18'b1000011000010111_00;
      patterns[1597] = 18'b1001011000010111_01;
      patterns[1598] = 18'b1010011000010111_10;
      patterns[1599] = 18'b1011011000010111_11;
      patterns[1600] = 18'b1000011000100000_00;
      patterns[1601] = 18'b1001011000100000_01;
      patterns[1602] = 18'b1010011000100000_10;
      patterns[1603] = 18'b1011011000100000_11;
      patterns[1604] = 18'b1000011000100001_00;
      patterns[1605] = 18'b1001011000100001_01;
      patterns[1606] = 18'b1010011000100001_10;
      patterns[1607] = 18'b1011011000100001_11;
      patterns[1608] = 18'b1000011000100010_00;
      patterns[1609] = 18'b1001011000100010_01;
      patterns[1610] = 18'b1010011000100010_10;
      patterns[1611] = 18'b1011011000100010_11;
      patterns[1612] = 18'b1000011000100011_00;
      patterns[1613] = 18'b1001011000100011_01;
      patterns[1614] = 18'b1010011000100011_10;
      patterns[1615] = 18'b1011011000100011_11;
      patterns[1616] = 18'b1000011000100100_00;
      patterns[1617] = 18'b1001011000100100_01;
      patterns[1618] = 18'b1010011000100100_10;
      patterns[1619] = 18'b1011011000100100_11;
      patterns[1620] = 18'b1000011000100101_00;
      patterns[1621] = 18'b1001011000100101_01;
      patterns[1622] = 18'b1010011000100101_10;
      patterns[1623] = 18'b1011011000100101_11;
      patterns[1624] = 18'b1000011000100110_00;
      patterns[1625] = 18'b1001011000100110_01;
      patterns[1626] = 18'b1010011000100110_10;
      patterns[1627] = 18'b1011011000100110_11;
      patterns[1628] = 18'b1000011000100111_00;
      patterns[1629] = 18'b1001011000100111_01;
      patterns[1630] = 18'b1010011000100111_10;
      patterns[1631] = 18'b1011011000100111_11;
      patterns[1632] = 18'b1000011000110000_00;
      patterns[1633] = 18'b1001011000110000_01;
      patterns[1634] = 18'b1010011000110000_10;
      patterns[1635] = 18'b1011011000110000_11;
      patterns[1636] = 18'b1000011000110001_00;
      patterns[1637] = 18'b1001011000110001_01;
      patterns[1638] = 18'b1010011000110001_10;
      patterns[1639] = 18'b1011011000110001_11;
      patterns[1640] = 18'b1000011000110010_00;
      patterns[1641] = 18'b1001011000110010_01;
      patterns[1642] = 18'b1010011000110010_10;
      patterns[1643] = 18'b1011011000110010_11;
      patterns[1644] = 18'b1000011000110011_00;
      patterns[1645] = 18'b1001011000110011_01;
      patterns[1646] = 18'b1010011000110011_10;
      patterns[1647] = 18'b1011011000110011_11;
      patterns[1648] = 18'b1000011000110100_00;
      patterns[1649] = 18'b1001011000110100_01;
      patterns[1650] = 18'b1010011000110100_10;
      patterns[1651] = 18'b1011011000110100_11;
      patterns[1652] = 18'b1000011000110101_00;
      patterns[1653] = 18'b1001011000110101_01;
      patterns[1654] = 18'b1010011000110101_10;
      patterns[1655] = 18'b1011011000110101_11;
      patterns[1656] = 18'b1000011000110110_00;
      patterns[1657] = 18'b1001011000110110_01;
      patterns[1658] = 18'b1010011000110110_10;
      patterns[1659] = 18'b1011011000110110_11;
      patterns[1660] = 18'b1000011000110111_00;
      patterns[1661] = 18'b1001011000110111_01;
      patterns[1662] = 18'b1010011000110111_10;
      patterns[1663] = 18'b1011011000110111_11;
      patterns[1664] = 18'b1000011001000000_00;
      patterns[1665] = 18'b1001011001000000_01;
      patterns[1666] = 18'b1010011001000000_10;
      patterns[1667] = 18'b1011011001000000_11;
      patterns[1668] = 18'b1000011001000001_00;
      patterns[1669] = 18'b1001011001000001_01;
      patterns[1670] = 18'b1010011001000001_10;
      patterns[1671] = 18'b1011011001000001_11;
      patterns[1672] = 18'b1000011001000010_00;
      patterns[1673] = 18'b1001011001000010_01;
      patterns[1674] = 18'b1010011001000010_10;
      patterns[1675] = 18'b1011011001000010_11;
      patterns[1676] = 18'b1000011001000011_00;
      patterns[1677] = 18'b1001011001000011_01;
      patterns[1678] = 18'b1010011001000011_10;
      patterns[1679] = 18'b1011011001000011_11;
      patterns[1680] = 18'b1000011001000100_00;
      patterns[1681] = 18'b1001011001000100_01;
      patterns[1682] = 18'b1010011001000100_10;
      patterns[1683] = 18'b1011011001000100_11;
      patterns[1684] = 18'b1000011001000101_00;
      patterns[1685] = 18'b1001011001000101_01;
      patterns[1686] = 18'b1010011001000101_10;
      patterns[1687] = 18'b1011011001000101_11;
      patterns[1688] = 18'b1000011001000110_00;
      patterns[1689] = 18'b1001011001000110_01;
      patterns[1690] = 18'b1010011001000110_10;
      patterns[1691] = 18'b1011011001000110_11;
      patterns[1692] = 18'b1000011001000111_00;
      patterns[1693] = 18'b1001011001000111_01;
      patterns[1694] = 18'b1010011001000111_10;
      patterns[1695] = 18'b1011011001000111_11;
      patterns[1696] = 18'b1000011001010000_00;
      patterns[1697] = 18'b1001011001010000_01;
      patterns[1698] = 18'b1010011001010000_10;
      patterns[1699] = 18'b1011011001010000_11;
      patterns[1700] = 18'b1000011001010001_00;
      patterns[1701] = 18'b1001011001010001_01;
      patterns[1702] = 18'b1010011001010001_10;
      patterns[1703] = 18'b1011011001010001_11;
      patterns[1704] = 18'b1000011001010010_00;
      patterns[1705] = 18'b1001011001010010_01;
      patterns[1706] = 18'b1010011001010010_10;
      patterns[1707] = 18'b1011011001010010_11;
      patterns[1708] = 18'b1000011001010011_00;
      patterns[1709] = 18'b1001011001010011_01;
      patterns[1710] = 18'b1010011001010011_10;
      patterns[1711] = 18'b1011011001010011_11;
      patterns[1712] = 18'b1000011001010100_00;
      patterns[1713] = 18'b1001011001010100_01;
      patterns[1714] = 18'b1010011001010100_10;
      patterns[1715] = 18'b1011011001010100_11;
      patterns[1716] = 18'b1000011001010101_00;
      patterns[1717] = 18'b1001011001010101_01;
      patterns[1718] = 18'b1010011001010101_10;
      patterns[1719] = 18'b1011011001010101_11;
      patterns[1720] = 18'b1000011001010110_00;
      patterns[1721] = 18'b1001011001010110_01;
      patterns[1722] = 18'b1010011001010110_10;
      patterns[1723] = 18'b1011011001010110_11;
      patterns[1724] = 18'b1000011001010111_00;
      patterns[1725] = 18'b1001011001010111_01;
      patterns[1726] = 18'b1010011001010111_10;
      patterns[1727] = 18'b1011011001010111_11;
      patterns[1728] = 18'b1000011001100000_00;
      patterns[1729] = 18'b1001011001100000_01;
      patterns[1730] = 18'b1010011001100000_10;
      patterns[1731] = 18'b1011011001100000_11;
      patterns[1732] = 18'b1000011001100001_00;
      patterns[1733] = 18'b1001011001100001_01;
      patterns[1734] = 18'b1010011001100001_10;
      patterns[1735] = 18'b1011011001100001_11;
      patterns[1736] = 18'b1000011001100010_00;
      patterns[1737] = 18'b1001011001100010_01;
      patterns[1738] = 18'b1010011001100010_10;
      patterns[1739] = 18'b1011011001100010_11;
      patterns[1740] = 18'b1000011001100011_00;
      patterns[1741] = 18'b1001011001100011_01;
      patterns[1742] = 18'b1010011001100011_10;
      patterns[1743] = 18'b1011011001100011_11;
      patterns[1744] = 18'b1000011001100100_00;
      patterns[1745] = 18'b1001011001100100_01;
      patterns[1746] = 18'b1010011001100100_10;
      patterns[1747] = 18'b1011011001100100_11;
      patterns[1748] = 18'b1000011001100101_00;
      patterns[1749] = 18'b1001011001100101_01;
      patterns[1750] = 18'b1010011001100101_10;
      patterns[1751] = 18'b1011011001100101_11;
      patterns[1752] = 18'b1000011001100110_00;
      patterns[1753] = 18'b1001011001100110_01;
      patterns[1754] = 18'b1010011001100110_10;
      patterns[1755] = 18'b1011011001100110_11;
      patterns[1756] = 18'b1000011001100111_00;
      patterns[1757] = 18'b1001011001100111_01;
      patterns[1758] = 18'b1010011001100111_10;
      patterns[1759] = 18'b1011011001100111_11;
      patterns[1760] = 18'b1000011001110000_00;
      patterns[1761] = 18'b1001011001110000_01;
      patterns[1762] = 18'b1010011001110000_10;
      patterns[1763] = 18'b1011011001110000_11;
      patterns[1764] = 18'b1000011001110001_00;
      patterns[1765] = 18'b1001011001110001_01;
      patterns[1766] = 18'b1010011001110001_10;
      patterns[1767] = 18'b1011011001110001_11;
      patterns[1768] = 18'b1000011001110010_00;
      patterns[1769] = 18'b1001011001110010_01;
      patterns[1770] = 18'b1010011001110010_10;
      patterns[1771] = 18'b1011011001110010_11;
      patterns[1772] = 18'b1000011001110011_00;
      patterns[1773] = 18'b1001011001110011_01;
      patterns[1774] = 18'b1010011001110011_10;
      patterns[1775] = 18'b1011011001110011_11;
      patterns[1776] = 18'b1000011001110100_00;
      patterns[1777] = 18'b1001011001110100_01;
      patterns[1778] = 18'b1010011001110100_10;
      patterns[1779] = 18'b1011011001110100_11;
      patterns[1780] = 18'b1000011001110101_00;
      patterns[1781] = 18'b1001011001110101_01;
      patterns[1782] = 18'b1010011001110101_10;
      patterns[1783] = 18'b1011011001110101_11;
      patterns[1784] = 18'b1000011001110110_00;
      patterns[1785] = 18'b1001011001110110_01;
      patterns[1786] = 18'b1010011001110110_10;
      patterns[1787] = 18'b1011011001110110_11;
      patterns[1788] = 18'b1000011001110111_00;
      patterns[1789] = 18'b1001011001110111_01;
      patterns[1790] = 18'b1010011001110111_10;
      patterns[1791] = 18'b1011011001110111_11;
      patterns[1792] = 18'b1000011100000000_00;
      patterns[1793] = 18'b1001011100000000_01;
      patterns[1794] = 18'b1010011100000000_10;
      patterns[1795] = 18'b1011011100000000_11;
      patterns[1796] = 18'b1000011100000001_00;
      patterns[1797] = 18'b1001011100000001_01;
      patterns[1798] = 18'b1010011100000001_10;
      patterns[1799] = 18'b1011011100000001_11;
      patterns[1800] = 18'b1000011100000010_00;
      patterns[1801] = 18'b1001011100000010_01;
      patterns[1802] = 18'b1010011100000010_10;
      patterns[1803] = 18'b1011011100000010_11;
      patterns[1804] = 18'b1000011100000011_00;
      patterns[1805] = 18'b1001011100000011_01;
      patterns[1806] = 18'b1010011100000011_10;
      patterns[1807] = 18'b1011011100000011_11;
      patterns[1808] = 18'b1000011100000100_00;
      patterns[1809] = 18'b1001011100000100_01;
      patterns[1810] = 18'b1010011100000100_10;
      patterns[1811] = 18'b1011011100000100_11;
      patterns[1812] = 18'b1000011100000101_00;
      patterns[1813] = 18'b1001011100000101_01;
      patterns[1814] = 18'b1010011100000101_10;
      patterns[1815] = 18'b1011011100000101_11;
      patterns[1816] = 18'b1000011100000110_00;
      patterns[1817] = 18'b1001011100000110_01;
      patterns[1818] = 18'b1010011100000110_10;
      patterns[1819] = 18'b1011011100000110_11;
      patterns[1820] = 18'b1000011100000111_00;
      patterns[1821] = 18'b1001011100000111_01;
      patterns[1822] = 18'b1010011100000111_10;
      patterns[1823] = 18'b1011011100000111_11;
      patterns[1824] = 18'b1000011100010000_00;
      patterns[1825] = 18'b1001011100010000_01;
      patterns[1826] = 18'b1010011100010000_10;
      patterns[1827] = 18'b1011011100010000_11;
      patterns[1828] = 18'b1000011100010001_00;
      patterns[1829] = 18'b1001011100010001_01;
      patterns[1830] = 18'b1010011100010001_10;
      patterns[1831] = 18'b1011011100010001_11;
      patterns[1832] = 18'b1000011100010010_00;
      patterns[1833] = 18'b1001011100010010_01;
      patterns[1834] = 18'b1010011100010010_10;
      patterns[1835] = 18'b1011011100010010_11;
      patterns[1836] = 18'b1000011100010011_00;
      patterns[1837] = 18'b1001011100010011_01;
      patterns[1838] = 18'b1010011100010011_10;
      patterns[1839] = 18'b1011011100010011_11;
      patterns[1840] = 18'b1000011100010100_00;
      patterns[1841] = 18'b1001011100010100_01;
      patterns[1842] = 18'b1010011100010100_10;
      patterns[1843] = 18'b1011011100010100_11;
      patterns[1844] = 18'b1000011100010101_00;
      patterns[1845] = 18'b1001011100010101_01;
      patterns[1846] = 18'b1010011100010101_10;
      patterns[1847] = 18'b1011011100010101_11;
      patterns[1848] = 18'b1000011100010110_00;
      patterns[1849] = 18'b1001011100010110_01;
      patterns[1850] = 18'b1010011100010110_10;
      patterns[1851] = 18'b1011011100010110_11;
      patterns[1852] = 18'b1000011100010111_00;
      patterns[1853] = 18'b1001011100010111_01;
      patterns[1854] = 18'b1010011100010111_10;
      patterns[1855] = 18'b1011011100010111_11;
      patterns[1856] = 18'b1000011100100000_00;
      patterns[1857] = 18'b1001011100100000_01;
      patterns[1858] = 18'b1010011100100000_10;
      patterns[1859] = 18'b1011011100100000_11;
      patterns[1860] = 18'b1000011100100001_00;
      patterns[1861] = 18'b1001011100100001_01;
      patterns[1862] = 18'b1010011100100001_10;
      patterns[1863] = 18'b1011011100100001_11;
      patterns[1864] = 18'b1000011100100010_00;
      patterns[1865] = 18'b1001011100100010_01;
      patterns[1866] = 18'b1010011100100010_10;
      patterns[1867] = 18'b1011011100100010_11;
      patterns[1868] = 18'b1000011100100011_00;
      patterns[1869] = 18'b1001011100100011_01;
      patterns[1870] = 18'b1010011100100011_10;
      patterns[1871] = 18'b1011011100100011_11;
      patterns[1872] = 18'b1000011100100100_00;
      patterns[1873] = 18'b1001011100100100_01;
      patterns[1874] = 18'b1010011100100100_10;
      patterns[1875] = 18'b1011011100100100_11;
      patterns[1876] = 18'b1000011100100101_00;
      patterns[1877] = 18'b1001011100100101_01;
      patterns[1878] = 18'b1010011100100101_10;
      patterns[1879] = 18'b1011011100100101_11;
      patterns[1880] = 18'b1000011100100110_00;
      patterns[1881] = 18'b1001011100100110_01;
      patterns[1882] = 18'b1010011100100110_10;
      patterns[1883] = 18'b1011011100100110_11;
      patterns[1884] = 18'b1000011100100111_00;
      patterns[1885] = 18'b1001011100100111_01;
      patterns[1886] = 18'b1010011100100111_10;
      patterns[1887] = 18'b1011011100100111_11;
      patterns[1888] = 18'b1000011100110000_00;
      patterns[1889] = 18'b1001011100110000_01;
      patterns[1890] = 18'b1010011100110000_10;
      patterns[1891] = 18'b1011011100110000_11;
      patterns[1892] = 18'b1000011100110001_00;
      patterns[1893] = 18'b1001011100110001_01;
      patterns[1894] = 18'b1010011100110001_10;
      patterns[1895] = 18'b1011011100110001_11;
      patterns[1896] = 18'b1000011100110010_00;
      patterns[1897] = 18'b1001011100110010_01;
      patterns[1898] = 18'b1010011100110010_10;
      patterns[1899] = 18'b1011011100110010_11;
      patterns[1900] = 18'b1000011100110011_00;
      patterns[1901] = 18'b1001011100110011_01;
      patterns[1902] = 18'b1010011100110011_10;
      patterns[1903] = 18'b1011011100110011_11;
      patterns[1904] = 18'b1000011100110100_00;
      patterns[1905] = 18'b1001011100110100_01;
      patterns[1906] = 18'b1010011100110100_10;
      patterns[1907] = 18'b1011011100110100_11;
      patterns[1908] = 18'b1000011100110101_00;
      patterns[1909] = 18'b1001011100110101_01;
      patterns[1910] = 18'b1010011100110101_10;
      patterns[1911] = 18'b1011011100110101_11;
      patterns[1912] = 18'b1000011100110110_00;
      patterns[1913] = 18'b1001011100110110_01;
      patterns[1914] = 18'b1010011100110110_10;
      patterns[1915] = 18'b1011011100110110_11;
      patterns[1916] = 18'b1000011100110111_00;
      patterns[1917] = 18'b1001011100110111_01;
      patterns[1918] = 18'b1010011100110111_10;
      patterns[1919] = 18'b1011011100110111_11;
      patterns[1920] = 18'b1000011101000000_00;
      patterns[1921] = 18'b1001011101000000_01;
      patterns[1922] = 18'b1010011101000000_10;
      patterns[1923] = 18'b1011011101000000_11;
      patterns[1924] = 18'b1000011101000001_00;
      patterns[1925] = 18'b1001011101000001_01;
      patterns[1926] = 18'b1010011101000001_10;
      patterns[1927] = 18'b1011011101000001_11;
      patterns[1928] = 18'b1000011101000010_00;
      patterns[1929] = 18'b1001011101000010_01;
      patterns[1930] = 18'b1010011101000010_10;
      patterns[1931] = 18'b1011011101000010_11;
      patterns[1932] = 18'b1000011101000011_00;
      patterns[1933] = 18'b1001011101000011_01;
      patterns[1934] = 18'b1010011101000011_10;
      patterns[1935] = 18'b1011011101000011_11;
      patterns[1936] = 18'b1000011101000100_00;
      patterns[1937] = 18'b1001011101000100_01;
      patterns[1938] = 18'b1010011101000100_10;
      patterns[1939] = 18'b1011011101000100_11;
      patterns[1940] = 18'b1000011101000101_00;
      patterns[1941] = 18'b1001011101000101_01;
      patterns[1942] = 18'b1010011101000101_10;
      patterns[1943] = 18'b1011011101000101_11;
      patterns[1944] = 18'b1000011101000110_00;
      patterns[1945] = 18'b1001011101000110_01;
      patterns[1946] = 18'b1010011101000110_10;
      patterns[1947] = 18'b1011011101000110_11;
      patterns[1948] = 18'b1000011101000111_00;
      patterns[1949] = 18'b1001011101000111_01;
      patterns[1950] = 18'b1010011101000111_10;
      patterns[1951] = 18'b1011011101000111_11;
      patterns[1952] = 18'b1000011101010000_00;
      patterns[1953] = 18'b1001011101010000_01;
      patterns[1954] = 18'b1010011101010000_10;
      patterns[1955] = 18'b1011011101010000_11;
      patterns[1956] = 18'b1000011101010001_00;
      patterns[1957] = 18'b1001011101010001_01;
      patterns[1958] = 18'b1010011101010001_10;
      patterns[1959] = 18'b1011011101010001_11;
      patterns[1960] = 18'b1000011101010010_00;
      patterns[1961] = 18'b1001011101010010_01;
      patterns[1962] = 18'b1010011101010010_10;
      patterns[1963] = 18'b1011011101010010_11;
      patterns[1964] = 18'b1000011101010011_00;
      patterns[1965] = 18'b1001011101010011_01;
      patterns[1966] = 18'b1010011101010011_10;
      patterns[1967] = 18'b1011011101010011_11;
      patterns[1968] = 18'b1000011101010100_00;
      patterns[1969] = 18'b1001011101010100_01;
      patterns[1970] = 18'b1010011101010100_10;
      patterns[1971] = 18'b1011011101010100_11;
      patterns[1972] = 18'b1000011101010101_00;
      patterns[1973] = 18'b1001011101010101_01;
      patterns[1974] = 18'b1010011101010101_10;
      patterns[1975] = 18'b1011011101010101_11;
      patterns[1976] = 18'b1000011101010110_00;
      patterns[1977] = 18'b1001011101010110_01;
      patterns[1978] = 18'b1010011101010110_10;
      patterns[1979] = 18'b1011011101010110_11;
      patterns[1980] = 18'b1000011101010111_00;
      patterns[1981] = 18'b1001011101010111_01;
      patterns[1982] = 18'b1010011101010111_10;
      patterns[1983] = 18'b1011011101010111_11;
      patterns[1984] = 18'b1000011101100000_00;
      patterns[1985] = 18'b1001011101100000_01;
      patterns[1986] = 18'b1010011101100000_10;
      patterns[1987] = 18'b1011011101100000_11;
      patterns[1988] = 18'b1000011101100001_00;
      patterns[1989] = 18'b1001011101100001_01;
      patterns[1990] = 18'b1010011101100001_10;
      patterns[1991] = 18'b1011011101100001_11;
      patterns[1992] = 18'b1000011101100010_00;
      patterns[1993] = 18'b1001011101100010_01;
      patterns[1994] = 18'b1010011101100010_10;
      patterns[1995] = 18'b1011011101100010_11;
      patterns[1996] = 18'b1000011101100011_00;
      patterns[1997] = 18'b1001011101100011_01;
      patterns[1998] = 18'b1010011101100011_10;
      patterns[1999] = 18'b1011011101100011_11;
      patterns[2000] = 18'b1000011101100100_00;
      patterns[2001] = 18'b1001011101100100_01;
      patterns[2002] = 18'b1010011101100100_10;
      patterns[2003] = 18'b1011011101100100_11;
      patterns[2004] = 18'b1000011101100101_00;
      patterns[2005] = 18'b1001011101100101_01;
      patterns[2006] = 18'b1010011101100101_10;
      patterns[2007] = 18'b1011011101100101_11;
      patterns[2008] = 18'b1000011101100110_00;
      patterns[2009] = 18'b1001011101100110_01;
      patterns[2010] = 18'b1010011101100110_10;
      patterns[2011] = 18'b1011011101100110_11;
      patterns[2012] = 18'b1000011101100111_00;
      patterns[2013] = 18'b1001011101100111_01;
      patterns[2014] = 18'b1010011101100111_10;
      patterns[2015] = 18'b1011011101100111_11;
      patterns[2016] = 18'b1000011101110000_00;
      patterns[2017] = 18'b1001011101110000_01;
      patterns[2018] = 18'b1010011101110000_10;
      patterns[2019] = 18'b1011011101110000_11;
      patterns[2020] = 18'b1000011101110001_00;
      patterns[2021] = 18'b1001011101110001_01;
      patterns[2022] = 18'b1010011101110001_10;
      patterns[2023] = 18'b1011011101110001_11;
      patterns[2024] = 18'b1000011101110010_00;
      patterns[2025] = 18'b1001011101110010_01;
      patterns[2026] = 18'b1010011101110010_10;
      patterns[2027] = 18'b1011011101110010_11;
      patterns[2028] = 18'b1000011101110011_00;
      patterns[2029] = 18'b1001011101110011_01;
      patterns[2030] = 18'b1010011101110011_10;
      patterns[2031] = 18'b1011011101110011_11;
      patterns[2032] = 18'b1000011101110100_00;
      patterns[2033] = 18'b1001011101110100_01;
      patterns[2034] = 18'b1010011101110100_10;
      patterns[2035] = 18'b1011011101110100_11;
      patterns[2036] = 18'b1000011101110101_00;
      patterns[2037] = 18'b1001011101110101_01;
      patterns[2038] = 18'b1010011101110101_10;
      patterns[2039] = 18'b1011011101110101_11;
      patterns[2040] = 18'b1000011101110110_00;
      patterns[2041] = 18'b1001011101110110_01;
      patterns[2042] = 18'b1010011101110110_10;
      patterns[2043] = 18'b1011011101110110_11;
      patterns[2044] = 18'b1000011101110111_00;
      patterns[2045] = 18'b1001011101110111_01;
      patterns[2046] = 18'b1010011101110111_10;
      patterns[2047] = 18'b1011011101110111_11;

      for (i = 0; i < 2048; i = i + 1)
      begin
        INST = patterns[i][17:2];
        #10;
        if (patterns[i][1:0] !== 2'hx)
        begin
          if (ALUOP !== patterns[i][1:0])
          begin
            $display("%d:ALUOP: (assertion error). Expected %h, found %h", i, patterns[i][1:0], ALUOP);
            $finish;
          end
        end
      end

      $display("All tests passed.");
    end
    endmodule
