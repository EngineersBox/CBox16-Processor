//  A testbench for control_unit_All Tests_tb
`timescale 1us/1ns

module control_unit_All Tests_tb;
    reg [15:0] INST;
    wire [1:0] ALUOP;
    wire [2:0] RS1;
    wire [2:0] RS2;
    wire [2:0] WS;
    wire STR;
    wire WE;
    wire [1:0] DMUX;
    wire LDR;

  control_unit control_unit0 (
    .INST(INST),
    .ALUOP(ALUOP),
    .RS1(RS1),
    .RS2(RS2),
    .WS(WS),
    .STR(STR),
    .WE(WE),
    .DMUX(DMUX),
    .LDR(LDR)
  );

    reg [31:0] patterns[0:3583];
    integer i;

    initial begin
      patterns[0] = 32'b1000000000000000_1_00_000_000_000_0_x_00;
      patterns[1] = 32'b1001000000000000_1_01_000_000_000_0_x_00;
      patterns[2] = 32'b1010000000000000_1_10_000_000_000_0_x_00;
      patterns[3] = 32'b1011000000000000_1_11_000_000_000_0_x_00;
      patterns[4] = 32'b0101000000000000_1_xx_000_xxx_000_0_1_01;
      patterns[5] = 32'b0100000000000000_0_xx_000_000_xxx_1_x_xx;
      patterns[6] = 32'b0000000001000010_1_xx_xxx_xxx_000_0_x_10;
      patterns[7] = 32'b1000000000000001_1_00_000_001_000_0_x_00;
      patterns[8] = 32'b1001000000000001_1_01_000_001_000_0_x_00;
      patterns[9] = 32'b1010000000000001_1_10_000_001_000_0_x_00;
      patterns[10] = 32'b1011000000000001_1_11_000_001_000_0_x_00;
      patterns[11] = 32'b0101000000000000_1_xx_000_xxx_000_0_1_01;
      patterns[12] = 32'b0100000000000000_0_xx_000_000_xxx_1_x_xx;
      patterns[13] = 32'b0000000001011101_1_xx_xxx_xxx_000_0_x_10;
      patterns[14] = 32'b1000000000000010_1_00_000_010_000_0_x_00;
      patterns[15] = 32'b1001000000000010_1_01_000_010_000_0_x_00;
      patterns[16] = 32'b1010000000000010_1_10_000_010_000_0_x_00;
      patterns[17] = 32'b1011000000000010_1_11_000_010_000_0_x_00;
      patterns[18] = 32'b0101000000000000_1_xx_000_xxx_000_0_1_01;
      patterns[19] = 32'b0100000000000000_0_xx_000_000_xxx_1_x_xx;
      patterns[20] = 32'b0000000011101010_1_xx_xxx_xxx_000_0_x_10;
      patterns[21] = 32'b1000000000000011_1_00_000_011_000_0_x_00;
      patterns[22] = 32'b1001000000000011_1_01_000_011_000_0_x_00;
      patterns[23] = 32'b1010000000000011_1_10_000_011_000_0_x_00;
      patterns[24] = 32'b1011000000000011_1_11_000_011_000_0_x_00;
      patterns[25] = 32'b0101000000000000_1_xx_000_xxx_000_0_1_01;
      patterns[26] = 32'b0100000000000000_0_xx_000_000_xxx_1_x_xx;
      patterns[27] = 32'b0000000010111101_1_xx_xxx_xxx_000_0_x_10;
      patterns[28] = 32'b1000000000000100_1_00_000_100_000_0_x_00;
      patterns[29] = 32'b1001000000000100_1_01_000_100_000_0_x_00;
      patterns[30] = 32'b1010000000000100_1_10_000_100_000_0_x_00;
      patterns[31] = 32'b1011000000000100_1_11_000_100_000_0_x_00;
      patterns[32] = 32'b0101000000000000_1_xx_000_xxx_000_0_1_01;
      patterns[33] = 32'b0100000000000000_0_xx_000_000_xxx_1_x_xx;
      patterns[34] = 32'b0000000010101101_1_xx_xxx_xxx_000_0_x_10;
      patterns[35] = 32'b1000000000000101_1_00_000_101_000_0_x_00;
      patterns[36] = 32'b1001000000000101_1_01_000_101_000_0_x_00;
      patterns[37] = 32'b1010000000000101_1_10_000_101_000_0_x_00;
      patterns[38] = 32'b1011000000000101_1_11_000_101_000_0_x_00;
      patterns[39] = 32'b0101000000000000_1_xx_000_xxx_000_0_1_01;
      patterns[40] = 32'b0100000000000000_0_xx_000_000_xxx_1_x_xx;
      patterns[41] = 32'b0000000010010110_1_xx_xxx_xxx_000_0_x_10;
      patterns[42] = 32'b1000000000000110_1_00_000_110_000_0_x_00;
      patterns[43] = 32'b1001000000000110_1_01_000_110_000_0_x_00;
      patterns[44] = 32'b1010000000000110_1_10_000_110_000_0_x_00;
      patterns[45] = 32'b1011000000000110_1_11_000_110_000_0_x_00;
      patterns[46] = 32'b0101000000000000_1_xx_000_xxx_000_0_1_01;
      patterns[47] = 32'b0100000000000000_0_xx_000_000_xxx_1_x_xx;
      patterns[48] = 32'b0000000011100101_1_xx_xxx_xxx_000_0_x_10;
      patterns[49] = 32'b1000000000000111_1_00_000_111_000_0_x_00;
      patterns[50] = 32'b1001000000000111_1_01_000_111_000_0_x_00;
      patterns[51] = 32'b1010000000000111_1_10_000_111_000_0_x_00;
      patterns[52] = 32'b1011000000000111_1_11_000_111_000_0_x_00;
      patterns[53] = 32'b0101000000000000_1_xx_000_xxx_000_0_1_01;
      patterns[54] = 32'b0100000000000000_0_xx_000_000_xxx_1_x_xx;
      patterns[55] = 32'b0000000001000011_1_xx_xxx_xxx_000_0_x_10;
      patterns[56] = 32'b1000000000010000_1_00_001_000_000_0_x_00;
      patterns[57] = 32'b1001000000010000_1_01_001_000_000_0_x_00;
      patterns[58] = 32'b1010000000010000_1_10_001_000_000_0_x_00;
      patterns[59] = 32'b1011000000010000_1_11_001_000_000_0_x_00;
      patterns[60] = 32'b0101000000010000_1_xx_001_xxx_000_0_1_01;
      patterns[61] = 32'b0100000000010000_0_xx_001_000_xxx_1_x_xx;
      patterns[62] = 32'b0000000000001100_1_xx_xxx_xxx_000_0_x_10;
      patterns[63] = 32'b1000000000010001_1_00_001_001_000_0_x_00;
      patterns[64] = 32'b1001000000010001_1_01_001_001_000_0_x_00;
      patterns[65] = 32'b1010000000010001_1_10_001_001_000_0_x_00;
      patterns[66] = 32'b1011000000010001_1_11_001_001_000_0_x_00;
      patterns[67] = 32'b0101000000010000_1_xx_001_xxx_000_0_1_01;
      patterns[68] = 32'b0100000000010000_0_xx_001_000_xxx_1_x_xx;
      patterns[69] = 32'b0000000010100001_1_xx_xxx_xxx_000_0_x_10;
      patterns[70] = 32'b1000000000010010_1_00_001_010_000_0_x_00;
      patterns[71] = 32'b1001000000010010_1_01_001_010_000_0_x_00;
      patterns[72] = 32'b1010000000010010_1_10_001_010_000_0_x_00;
      patterns[73] = 32'b1011000000010010_1_11_001_010_000_0_x_00;
      patterns[74] = 32'b0101000000010000_1_xx_001_xxx_000_0_1_01;
      patterns[75] = 32'b0100000000010000_0_xx_001_000_xxx_1_x_xx;
      patterns[76] = 32'b0000000000011111_1_xx_xxx_xxx_000_0_x_10;
      patterns[77] = 32'b1000000000010011_1_00_001_011_000_0_x_00;
      patterns[78] = 32'b1001000000010011_1_01_001_011_000_0_x_00;
      patterns[79] = 32'b1010000000010011_1_10_001_011_000_0_x_00;
      patterns[80] = 32'b1011000000010011_1_11_001_011_000_0_x_00;
      patterns[81] = 32'b0101000000010000_1_xx_001_xxx_000_0_1_01;
      patterns[82] = 32'b0100000000010000_0_xx_001_000_xxx_1_x_xx;
      patterns[83] = 32'b0000000011110111_1_xx_xxx_xxx_000_0_x_10;
      patterns[84] = 32'b1000000000010100_1_00_001_100_000_0_x_00;
      patterns[85] = 32'b1001000000010100_1_01_001_100_000_0_x_00;
      patterns[86] = 32'b1010000000010100_1_10_001_100_000_0_x_00;
      patterns[87] = 32'b1011000000010100_1_11_001_100_000_0_x_00;
      patterns[88] = 32'b0101000000010000_1_xx_001_xxx_000_0_1_01;
      patterns[89] = 32'b0100000000010000_0_xx_001_000_xxx_1_x_xx;
      patterns[90] = 32'b0000000011100110_1_xx_xxx_xxx_000_0_x_10;
      patterns[91] = 32'b1000000000010101_1_00_001_101_000_0_x_00;
      patterns[92] = 32'b1001000000010101_1_01_001_101_000_0_x_00;
      patterns[93] = 32'b1010000000010101_1_10_001_101_000_0_x_00;
      patterns[94] = 32'b1011000000010101_1_11_001_101_000_0_x_00;
      patterns[95] = 32'b0101000000010000_1_xx_001_xxx_000_0_1_01;
      patterns[96] = 32'b0100000000010000_0_xx_001_000_xxx_1_x_xx;
      patterns[97] = 32'b0000000000001111_1_xx_xxx_xxx_000_0_x_10;
      patterns[98] = 32'b1000000000010110_1_00_001_110_000_0_x_00;
      patterns[99] = 32'b1001000000010110_1_01_001_110_000_0_x_00;
      patterns[100] = 32'b1010000000010110_1_10_001_110_000_0_x_00;
      patterns[101] = 32'b1011000000010110_1_11_001_110_000_0_x_00;
      patterns[102] = 32'b0101000000010000_1_xx_001_xxx_000_0_1_01;
      patterns[103] = 32'b0100000000010000_0_xx_001_000_xxx_1_x_xx;
      patterns[104] = 32'b0000000000000000_1_xx_xxx_xxx_000_0_x_10;
      patterns[105] = 32'b1000000000010111_1_00_001_111_000_0_x_00;
      patterns[106] = 32'b1001000000010111_1_01_001_111_000_0_x_00;
      patterns[107] = 32'b1010000000010111_1_10_001_111_000_0_x_00;
      patterns[108] = 32'b1011000000010111_1_11_001_111_000_0_x_00;
      patterns[109] = 32'b0101000000010000_1_xx_001_xxx_000_0_1_01;
      patterns[110] = 32'b0100000000010000_0_xx_001_000_xxx_1_x_xx;
      patterns[111] = 32'b0000000001011000_1_xx_xxx_xxx_000_0_x_10;
      patterns[112] = 32'b1000000000100000_1_00_010_000_000_0_x_00;
      patterns[113] = 32'b1001000000100000_1_01_010_000_000_0_x_00;
      patterns[114] = 32'b1010000000100000_1_10_010_000_000_0_x_00;
      patterns[115] = 32'b1011000000100000_1_11_010_000_000_0_x_00;
      patterns[116] = 32'b0101000000100000_1_xx_010_xxx_000_0_1_01;
      patterns[117] = 32'b0100000000100000_0_xx_010_000_xxx_1_x_xx;
      patterns[118] = 32'b0000000001011000_1_xx_xxx_xxx_000_0_x_10;
      patterns[119] = 32'b1000000000100001_1_00_010_001_000_0_x_00;
      patterns[120] = 32'b1001000000100001_1_01_010_001_000_0_x_00;
      patterns[121] = 32'b1010000000100001_1_10_010_001_000_0_x_00;
      patterns[122] = 32'b1011000000100001_1_11_010_001_000_0_x_00;
      patterns[123] = 32'b0101000000100000_1_xx_010_xxx_000_0_1_01;
      patterns[124] = 32'b0100000000100000_0_xx_010_000_xxx_1_x_xx;
      patterns[125] = 32'b0000000010001011_1_xx_xxx_xxx_000_0_x_10;
      patterns[126] = 32'b1000000000100010_1_00_010_010_000_0_x_00;
      patterns[127] = 32'b1001000000100010_1_01_010_010_000_0_x_00;
      patterns[128] = 32'b1010000000100010_1_10_010_010_000_0_x_00;
      patterns[129] = 32'b1011000000100010_1_11_010_010_000_0_x_00;
      patterns[130] = 32'b0101000000100000_1_xx_010_xxx_000_0_1_01;
      patterns[131] = 32'b0100000000100000_0_xx_010_000_xxx_1_x_xx;
      patterns[132] = 32'b0000000001000111_1_xx_xxx_xxx_000_0_x_10;
      patterns[133] = 32'b1000000000100011_1_00_010_011_000_0_x_00;
      patterns[134] = 32'b1001000000100011_1_01_010_011_000_0_x_00;
      patterns[135] = 32'b1010000000100011_1_10_010_011_000_0_x_00;
      patterns[136] = 32'b1011000000100011_1_11_010_011_000_0_x_00;
      patterns[137] = 32'b0101000000100000_1_xx_010_xxx_000_0_1_01;
      patterns[138] = 32'b0100000000100000_0_xx_010_000_xxx_1_x_xx;
      patterns[139] = 32'b0000000000100100_1_xx_xxx_xxx_000_0_x_10;
      patterns[140] = 32'b1000000000100100_1_00_010_100_000_0_x_00;
      patterns[141] = 32'b1001000000100100_1_01_010_100_000_0_x_00;
      patterns[142] = 32'b1010000000100100_1_10_010_100_000_0_x_00;
      patterns[143] = 32'b1011000000100100_1_11_010_100_000_0_x_00;
      patterns[144] = 32'b0101000000100000_1_xx_010_xxx_000_0_1_01;
      patterns[145] = 32'b0100000000100000_0_xx_010_000_xxx_1_x_xx;
      patterns[146] = 32'b0000000011101001_1_xx_xxx_xxx_000_0_x_10;
      patterns[147] = 32'b1000000000100101_1_00_010_101_000_0_x_00;
      patterns[148] = 32'b1001000000100101_1_01_010_101_000_0_x_00;
      patterns[149] = 32'b1010000000100101_1_10_010_101_000_0_x_00;
      patterns[150] = 32'b1011000000100101_1_11_010_101_000_0_x_00;
      patterns[151] = 32'b0101000000100000_1_xx_010_xxx_000_0_1_01;
      patterns[152] = 32'b0100000000100000_0_xx_010_000_xxx_1_x_xx;
      patterns[153] = 32'b0000000001100000_1_xx_xxx_xxx_000_0_x_10;
      patterns[154] = 32'b1000000000100110_1_00_010_110_000_0_x_00;
      patterns[155] = 32'b1001000000100110_1_01_010_110_000_0_x_00;
      patterns[156] = 32'b1010000000100110_1_10_010_110_000_0_x_00;
      patterns[157] = 32'b1011000000100110_1_11_010_110_000_0_x_00;
      patterns[158] = 32'b0101000000100000_1_xx_010_xxx_000_0_1_01;
      patterns[159] = 32'b0100000000100000_0_xx_010_000_xxx_1_x_xx;
      patterns[160] = 32'b0000000001001100_1_xx_xxx_xxx_000_0_x_10;
      patterns[161] = 32'b1000000000100111_1_00_010_111_000_0_x_00;
      patterns[162] = 32'b1001000000100111_1_01_010_111_000_0_x_00;
      patterns[163] = 32'b1010000000100111_1_10_010_111_000_0_x_00;
      patterns[164] = 32'b1011000000100111_1_11_010_111_000_0_x_00;
      patterns[165] = 32'b0101000000100000_1_xx_010_xxx_000_0_1_01;
      patterns[166] = 32'b0100000000100000_0_xx_010_000_xxx_1_x_xx;
      patterns[167] = 32'b0000000010110000_1_xx_xxx_xxx_000_0_x_10;
      patterns[168] = 32'b1000000000110000_1_00_011_000_000_0_x_00;
      patterns[169] = 32'b1001000000110000_1_01_011_000_000_0_x_00;
      patterns[170] = 32'b1010000000110000_1_10_011_000_000_0_x_00;
      patterns[171] = 32'b1011000000110000_1_11_011_000_000_0_x_00;
      patterns[172] = 32'b0101000000110000_1_xx_011_xxx_000_0_1_01;
      patterns[173] = 32'b0100000000110000_0_xx_011_000_xxx_1_x_xx;
      patterns[174] = 32'b0000000000000111_1_xx_xxx_xxx_000_0_x_10;
      patterns[175] = 32'b1000000000110001_1_00_011_001_000_0_x_00;
      patterns[176] = 32'b1001000000110001_1_01_011_001_000_0_x_00;
      patterns[177] = 32'b1010000000110001_1_10_011_001_000_0_x_00;
      patterns[178] = 32'b1011000000110001_1_11_011_001_000_0_x_00;
      patterns[179] = 32'b0101000000110000_1_xx_011_xxx_000_0_1_01;
      patterns[180] = 32'b0100000000110000_0_xx_011_000_xxx_1_x_xx;
      patterns[181] = 32'b0000000011010110_1_xx_xxx_xxx_000_0_x_10;
      patterns[182] = 32'b1000000000110010_1_00_011_010_000_0_x_00;
      patterns[183] = 32'b1001000000110010_1_01_011_010_000_0_x_00;
      patterns[184] = 32'b1010000000110010_1_10_011_010_000_0_x_00;
      patterns[185] = 32'b1011000000110010_1_11_011_010_000_0_x_00;
      patterns[186] = 32'b0101000000110000_1_xx_011_xxx_000_0_1_01;
      patterns[187] = 32'b0100000000110000_0_xx_011_000_xxx_1_x_xx;
      patterns[188] = 32'b0000000010101010_1_xx_xxx_xxx_000_0_x_10;
      patterns[189] = 32'b1000000000110011_1_00_011_011_000_0_x_00;
      patterns[190] = 32'b1001000000110011_1_01_011_011_000_0_x_00;
      patterns[191] = 32'b1010000000110011_1_10_011_011_000_0_x_00;
      patterns[192] = 32'b1011000000110011_1_11_011_011_000_0_x_00;
      patterns[193] = 32'b0101000000110000_1_xx_011_xxx_000_0_1_01;
      patterns[194] = 32'b0100000000110000_0_xx_011_000_xxx_1_x_xx;
      patterns[195] = 32'b0000000000000110_1_xx_xxx_xxx_000_0_x_10;
      patterns[196] = 32'b1000000000110100_1_00_011_100_000_0_x_00;
      patterns[197] = 32'b1001000000110100_1_01_011_100_000_0_x_00;
      patterns[198] = 32'b1010000000110100_1_10_011_100_000_0_x_00;
      patterns[199] = 32'b1011000000110100_1_11_011_100_000_0_x_00;
      patterns[200] = 32'b0101000000110000_1_xx_011_xxx_000_0_1_01;
      patterns[201] = 32'b0100000000110000_0_xx_011_000_xxx_1_x_xx;
      patterns[202] = 32'b0000000000100100_1_xx_xxx_xxx_000_0_x_10;
      patterns[203] = 32'b1000000000110101_1_00_011_101_000_0_x_00;
      patterns[204] = 32'b1001000000110101_1_01_011_101_000_0_x_00;
      patterns[205] = 32'b1010000000110101_1_10_011_101_000_0_x_00;
      patterns[206] = 32'b1011000000110101_1_11_011_101_000_0_x_00;
      patterns[207] = 32'b0101000000110000_1_xx_011_xxx_000_0_1_01;
      patterns[208] = 32'b0100000000110000_0_xx_011_000_xxx_1_x_xx;
      patterns[209] = 32'b0000000000110101_1_xx_xxx_xxx_000_0_x_10;
      patterns[210] = 32'b1000000000110110_1_00_011_110_000_0_x_00;
      patterns[211] = 32'b1001000000110110_1_01_011_110_000_0_x_00;
      patterns[212] = 32'b1010000000110110_1_10_011_110_000_0_x_00;
      patterns[213] = 32'b1011000000110110_1_11_011_110_000_0_x_00;
      patterns[214] = 32'b0101000000110000_1_xx_011_xxx_000_0_1_01;
      patterns[215] = 32'b0100000000110000_0_xx_011_000_xxx_1_x_xx;
      patterns[216] = 32'b0000000010000101_1_xx_xxx_xxx_000_0_x_10;
      patterns[217] = 32'b1000000000110111_1_00_011_111_000_0_x_00;
      patterns[218] = 32'b1001000000110111_1_01_011_111_000_0_x_00;
      patterns[219] = 32'b1010000000110111_1_10_011_111_000_0_x_00;
      patterns[220] = 32'b1011000000110111_1_11_011_111_000_0_x_00;
      patterns[221] = 32'b0101000000110000_1_xx_011_xxx_000_0_1_01;
      patterns[222] = 32'b0100000000110000_0_xx_011_000_xxx_1_x_xx;
      patterns[223] = 32'b0000000000001100_1_xx_xxx_xxx_000_0_x_10;
      patterns[224] = 32'b1000000001000000_1_00_100_000_000_0_x_00;
      patterns[225] = 32'b1001000001000000_1_01_100_000_000_0_x_00;
      patterns[226] = 32'b1010000001000000_1_10_100_000_000_0_x_00;
      patterns[227] = 32'b1011000001000000_1_11_100_000_000_0_x_00;
      patterns[228] = 32'b0101000001000000_1_xx_100_xxx_000_0_1_01;
      patterns[229] = 32'b0100000001000000_0_xx_100_000_xxx_1_x_xx;
      patterns[230] = 32'b0000000010001100_1_xx_xxx_xxx_000_0_x_10;
      patterns[231] = 32'b1000000001000001_1_00_100_001_000_0_x_00;
      patterns[232] = 32'b1001000001000001_1_01_100_001_000_0_x_00;
      patterns[233] = 32'b1010000001000001_1_10_100_001_000_0_x_00;
      patterns[234] = 32'b1011000001000001_1_11_100_001_000_0_x_00;
      patterns[235] = 32'b0101000001000000_1_xx_100_xxx_000_0_1_01;
      patterns[236] = 32'b0100000001000000_0_xx_100_000_xxx_1_x_xx;
      patterns[237] = 32'b0000000010011001_1_xx_xxx_xxx_000_0_x_10;
      patterns[238] = 32'b1000000001000010_1_00_100_010_000_0_x_00;
      patterns[239] = 32'b1001000001000010_1_01_100_010_000_0_x_00;
      patterns[240] = 32'b1010000001000010_1_10_100_010_000_0_x_00;
      patterns[241] = 32'b1011000001000010_1_11_100_010_000_0_x_00;
      patterns[242] = 32'b0101000001000000_1_xx_100_xxx_000_0_1_01;
      patterns[243] = 32'b0100000001000000_0_xx_100_000_xxx_1_x_xx;
      patterns[244] = 32'b0000000010100111_1_xx_xxx_xxx_000_0_x_10;
      patterns[245] = 32'b1000000001000011_1_00_100_011_000_0_x_00;
      patterns[246] = 32'b1001000001000011_1_01_100_011_000_0_x_00;
      patterns[247] = 32'b1010000001000011_1_10_100_011_000_0_x_00;
      patterns[248] = 32'b1011000001000011_1_11_100_011_000_0_x_00;
      patterns[249] = 32'b0101000001000000_1_xx_100_xxx_000_0_1_01;
      patterns[250] = 32'b0100000001000000_0_xx_100_000_xxx_1_x_xx;
      patterns[251] = 32'b0000000011110010_1_xx_xxx_xxx_000_0_x_10;
      patterns[252] = 32'b1000000001000100_1_00_100_100_000_0_x_00;
      patterns[253] = 32'b1001000001000100_1_01_100_100_000_0_x_00;
      patterns[254] = 32'b1010000001000100_1_10_100_100_000_0_x_00;
      patterns[255] = 32'b1011000001000100_1_11_100_100_000_0_x_00;
      patterns[256] = 32'b0101000001000000_1_xx_100_xxx_000_0_1_01;
      patterns[257] = 32'b0100000001000000_0_xx_100_000_xxx_1_x_xx;
      patterns[258] = 32'b0000000010110000_1_xx_xxx_xxx_000_0_x_10;
      patterns[259] = 32'b1000000001000101_1_00_100_101_000_0_x_00;
      patterns[260] = 32'b1001000001000101_1_01_100_101_000_0_x_00;
      patterns[261] = 32'b1010000001000101_1_10_100_101_000_0_x_00;
      patterns[262] = 32'b1011000001000101_1_11_100_101_000_0_x_00;
      patterns[263] = 32'b0101000001000000_1_xx_100_xxx_000_0_1_01;
      patterns[264] = 32'b0100000001000000_0_xx_100_000_xxx_1_x_xx;
      patterns[265] = 32'b0000000010101000_1_xx_xxx_xxx_000_0_x_10;
      patterns[266] = 32'b1000000001000110_1_00_100_110_000_0_x_00;
      patterns[267] = 32'b1001000001000110_1_01_100_110_000_0_x_00;
      patterns[268] = 32'b1010000001000110_1_10_100_110_000_0_x_00;
      patterns[269] = 32'b1011000001000110_1_11_100_110_000_0_x_00;
      patterns[270] = 32'b0101000001000000_1_xx_100_xxx_000_0_1_01;
      patterns[271] = 32'b0100000001000000_0_xx_100_000_xxx_1_x_xx;
      patterns[272] = 32'b0000000011010010_1_xx_xxx_xxx_000_0_x_10;
      patterns[273] = 32'b1000000001000111_1_00_100_111_000_0_x_00;
      patterns[274] = 32'b1001000001000111_1_01_100_111_000_0_x_00;
      patterns[275] = 32'b1010000001000111_1_10_100_111_000_0_x_00;
      patterns[276] = 32'b1011000001000111_1_11_100_111_000_0_x_00;
      patterns[277] = 32'b0101000001000000_1_xx_100_xxx_000_0_1_01;
      patterns[278] = 32'b0100000001000000_0_xx_100_000_xxx_1_x_xx;
      patterns[279] = 32'b0000000011111100_1_xx_xxx_xxx_000_0_x_10;
      patterns[280] = 32'b1000000001010000_1_00_101_000_000_0_x_00;
      patterns[281] = 32'b1001000001010000_1_01_101_000_000_0_x_00;
      patterns[282] = 32'b1010000001010000_1_10_101_000_000_0_x_00;
      patterns[283] = 32'b1011000001010000_1_11_101_000_000_0_x_00;
      patterns[284] = 32'b0101000001010000_1_xx_101_xxx_000_0_1_01;
      patterns[285] = 32'b0100000001010000_0_xx_101_000_xxx_1_x_xx;
      patterns[286] = 32'b0000000000010110_1_xx_xxx_xxx_000_0_x_10;
      patterns[287] = 32'b1000000001010001_1_00_101_001_000_0_x_00;
      patterns[288] = 32'b1001000001010001_1_01_101_001_000_0_x_00;
      patterns[289] = 32'b1010000001010001_1_10_101_001_000_0_x_00;
      patterns[290] = 32'b1011000001010001_1_11_101_001_000_0_x_00;
      patterns[291] = 32'b0101000001010000_1_xx_101_xxx_000_0_1_01;
      patterns[292] = 32'b0100000001010000_0_xx_101_000_xxx_1_x_xx;
      patterns[293] = 32'b0000000000110111_1_xx_xxx_xxx_000_0_x_10;
      patterns[294] = 32'b1000000001010010_1_00_101_010_000_0_x_00;
      patterns[295] = 32'b1001000001010010_1_01_101_010_000_0_x_00;
      patterns[296] = 32'b1010000001010010_1_10_101_010_000_0_x_00;
      patterns[297] = 32'b1011000001010010_1_11_101_010_000_0_x_00;
      patterns[298] = 32'b0101000001010000_1_xx_101_xxx_000_0_1_01;
      patterns[299] = 32'b0100000001010000_0_xx_101_000_xxx_1_x_xx;
      patterns[300] = 32'b0000000011101011_1_xx_xxx_xxx_000_0_x_10;
      patterns[301] = 32'b1000000001010011_1_00_101_011_000_0_x_00;
      patterns[302] = 32'b1001000001010011_1_01_101_011_000_0_x_00;
      patterns[303] = 32'b1010000001010011_1_10_101_011_000_0_x_00;
      patterns[304] = 32'b1011000001010011_1_11_101_011_000_0_x_00;
      patterns[305] = 32'b0101000001010000_1_xx_101_xxx_000_0_1_01;
      patterns[306] = 32'b0100000001010000_0_xx_101_000_xxx_1_x_xx;
      patterns[307] = 32'b0000000001110100_1_xx_xxx_xxx_000_0_x_10;
      patterns[308] = 32'b1000000001010100_1_00_101_100_000_0_x_00;
      patterns[309] = 32'b1001000001010100_1_01_101_100_000_0_x_00;
      patterns[310] = 32'b1010000001010100_1_10_101_100_000_0_x_00;
      patterns[311] = 32'b1011000001010100_1_11_101_100_000_0_x_00;
      patterns[312] = 32'b0101000001010000_1_xx_101_xxx_000_0_1_01;
      patterns[313] = 32'b0100000001010000_0_xx_101_000_xxx_1_x_xx;
      patterns[314] = 32'b0000000011110101_1_xx_xxx_xxx_000_0_x_10;
      patterns[315] = 32'b1000000001010101_1_00_101_101_000_0_x_00;
      patterns[316] = 32'b1001000001010101_1_01_101_101_000_0_x_00;
      patterns[317] = 32'b1010000001010101_1_10_101_101_000_0_x_00;
      patterns[318] = 32'b1011000001010101_1_11_101_101_000_0_x_00;
      patterns[319] = 32'b0101000001010000_1_xx_101_xxx_000_0_1_01;
      patterns[320] = 32'b0100000001010000_0_xx_101_000_xxx_1_x_xx;
      patterns[321] = 32'b0000000010101100_1_xx_xxx_xxx_000_0_x_10;
      patterns[322] = 32'b1000000001010110_1_00_101_110_000_0_x_00;
      patterns[323] = 32'b1001000001010110_1_01_101_110_000_0_x_00;
      patterns[324] = 32'b1010000001010110_1_10_101_110_000_0_x_00;
      patterns[325] = 32'b1011000001010110_1_11_101_110_000_0_x_00;
      patterns[326] = 32'b0101000001010000_1_xx_101_xxx_000_0_1_01;
      patterns[327] = 32'b0100000001010000_0_xx_101_000_xxx_1_x_xx;
      patterns[328] = 32'b0000000000101101_1_xx_xxx_xxx_000_0_x_10;
      patterns[329] = 32'b1000000001010111_1_00_101_111_000_0_x_00;
      patterns[330] = 32'b1001000001010111_1_01_101_111_000_0_x_00;
      patterns[331] = 32'b1010000001010111_1_10_101_111_000_0_x_00;
      patterns[332] = 32'b1011000001010111_1_11_101_111_000_0_x_00;
      patterns[333] = 32'b0101000001010000_1_xx_101_xxx_000_0_1_01;
      patterns[334] = 32'b0100000001010000_0_xx_101_000_xxx_1_x_xx;
      patterns[335] = 32'b0000000001001010_1_xx_xxx_xxx_000_0_x_10;
      patterns[336] = 32'b1000000001100000_1_00_110_000_000_0_x_00;
      patterns[337] = 32'b1001000001100000_1_01_110_000_000_0_x_00;
      patterns[338] = 32'b1010000001100000_1_10_110_000_000_0_x_00;
      patterns[339] = 32'b1011000001100000_1_11_110_000_000_0_x_00;
      patterns[340] = 32'b0101000001100000_1_xx_110_xxx_000_0_1_01;
      patterns[341] = 32'b0100000001100000_0_xx_110_000_xxx_1_x_xx;
      patterns[342] = 32'b0000000001101100_1_xx_xxx_xxx_000_0_x_10;
      patterns[343] = 32'b1000000001100001_1_00_110_001_000_0_x_00;
      patterns[344] = 32'b1001000001100001_1_01_110_001_000_0_x_00;
      patterns[345] = 32'b1010000001100001_1_10_110_001_000_0_x_00;
      patterns[346] = 32'b1011000001100001_1_11_110_001_000_0_x_00;
      patterns[347] = 32'b0101000001100000_1_xx_110_xxx_000_0_1_01;
      patterns[348] = 32'b0100000001100000_0_xx_110_000_xxx_1_x_xx;
      patterns[349] = 32'b0000000011001100_1_xx_xxx_xxx_000_0_x_10;
      patterns[350] = 32'b1000000001100010_1_00_110_010_000_0_x_00;
      patterns[351] = 32'b1001000001100010_1_01_110_010_000_0_x_00;
      patterns[352] = 32'b1010000001100010_1_10_110_010_000_0_x_00;
      patterns[353] = 32'b1011000001100010_1_11_110_010_000_0_x_00;
      patterns[354] = 32'b0101000001100000_1_xx_110_xxx_000_0_1_01;
      patterns[355] = 32'b0100000001100000_0_xx_110_000_xxx_1_x_xx;
      patterns[356] = 32'b0000000000010100_1_xx_xxx_xxx_000_0_x_10;
      patterns[357] = 32'b1000000001100011_1_00_110_011_000_0_x_00;
      patterns[358] = 32'b1001000001100011_1_01_110_011_000_0_x_00;
      patterns[359] = 32'b1010000001100011_1_10_110_011_000_0_x_00;
      patterns[360] = 32'b1011000001100011_1_11_110_011_000_0_x_00;
      patterns[361] = 32'b0101000001100000_1_xx_110_xxx_000_0_1_01;
      patterns[362] = 32'b0100000001100000_0_xx_110_000_xxx_1_x_xx;
      patterns[363] = 32'b0000000001101100_1_xx_xxx_xxx_000_0_x_10;
      patterns[364] = 32'b1000000001100100_1_00_110_100_000_0_x_00;
      patterns[365] = 32'b1001000001100100_1_01_110_100_000_0_x_00;
      patterns[366] = 32'b1010000001100100_1_10_110_100_000_0_x_00;
      patterns[367] = 32'b1011000001100100_1_11_110_100_000_0_x_00;
      patterns[368] = 32'b0101000001100000_1_xx_110_xxx_000_0_1_01;
      patterns[369] = 32'b0100000001100000_0_xx_110_000_xxx_1_x_xx;
      patterns[370] = 32'b0000000001010101_1_xx_xxx_xxx_000_0_x_10;
      patterns[371] = 32'b1000000001100101_1_00_110_101_000_0_x_00;
      patterns[372] = 32'b1001000001100101_1_01_110_101_000_0_x_00;
      patterns[373] = 32'b1010000001100101_1_10_110_101_000_0_x_00;
      patterns[374] = 32'b1011000001100101_1_11_110_101_000_0_x_00;
      patterns[375] = 32'b0101000001100000_1_xx_110_xxx_000_0_1_01;
      patterns[376] = 32'b0100000001100000_0_xx_110_000_xxx_1_x_xx;
      patterns[377] = 32'b0000000000010111_1_xx_xxx_xxx_000_0_x_10;
      patterns[378] = 32'b1000000001100110_1_00_110_110_000_0_x_00;
      patterns[379] = 32'b1001000001100110_1_01_110_110_000_0_x_00;
      patterns[380] = 32'b1010000001100110_1_10_110_110_000_0_x_00;
      patterns[381] = 32'b1011000001100110_1_11_110_110_000_0_x_00;
      patterns[382] = 32'b0101000001100000_1_xx_110_xxx_000_0_1_01;
      patterns[383] = 32'b0100000001100000_0_xx_110_000_xxx_1_x_xx;
      patterns[384] = 32'b0000000010100111_1_xx_xxx_xxx_000_0_x_10;
      patterns[385] = 32'b1000000001100111_1_00_110_111_000_0_x_00;
      patterns[386] = 32'b1001000001100111_1_01_110_111_000_0_x_00;
      patterns[387] = 32'b1010000001100111_1_10_110_111_000_0_x_00;
      patterns[388] = 32'b1011000001100111_1_11_110_111_000_0_x_00;
      patterns[389] = 32'b0101000001100000_1_xx_110_xxx_000_0_1_01;
      patterns[390] = 32'b0100000001100000_0_xx_110_000_xxx_1_x_xx;
      patterns[391] = 32'b0000000001011111_1_xx_xxx_xxx_000_0_x_10;
      patterns[392] = 32'b1000000001110000_1_00_111_000_000_0_x_00;
      patterns[393] = 32'b1001000001110000_1_01_111_000_000_0_x_00;
      patterns[394] = 32'b1010000001110000_1_10_111_000_000_0_x_00;
      patterns[395] = 32'b1011000001110000_1_11_111_000_000_0_x_00;
      patterns[396] = 32'b0101000001110000_1_xx_111_xxx_000_0_1_01;
      patterns[397] = 32'b0100000001110000_0_xx_111_000_xxx_1_x_xx;
      patterns[398] = 32'b0000000011101111_1_xx_xxx_xxx_000_0_x_10;
      patterns[399] = 32'b1000000001110001_1_00_111_001_000_0_x_00;
      patterns[400] = 32'b1001000001110001_1_01_111_001_000_0_x_00;
      patterns[401] = 32'b1010000001110001_1_10_111_001_000_0_x_00;
      patterns[402] = 32'b1011000001110001_1_11_111_001_000_0_x_00;
      patterns[403] = 32'b0101000001110000_1_xx_111_xxx_000_0_1_01;
      patterns[404] = 32'b0100000001110000_0_xx_111_000_xxx_1_x_xx;
      patterns[405] = 32'b0000000010011011_1_xx_xxx_xxx_000_0_x_10;
      patterns[406] = 32'b1000000001110010_1_00_111_010_000_0_x_00;
      patterns[407] = 32'b1001000001110010_1_01_111_010_000_0_x_00;
      patterns[408] = 32'b1010000001110010_1_10_111_010_000_0_x_00;
      patterns[409] = 32'b1011000001110010_1_11_111_010_000_0_x_00;
      patterns[410] = 32'b0101000001110000_1_xx_111_xxx_000_0_1_01;
      patterns[411] = 32'b0100000001110000_0_xx_111_000_xxx_1_x_xx;
      patterns[412] = 32'b0000000001111000_1_xx_xxx_xxx_000_0_x_10;
      patterns[413] = 32'b1000000001110011_1_00_111_011_000_0_x_00;
      patterns[414] = 32'b1001000001110011_1_01_111_011_000_0_x_00;
      patterns[415] = 32'b1010000001110011_1_10_111_011_000_0_x_00;
      patterns[416] = 32'b1011000001110011_1_11_111_011_000_0_x_00;
      patterns[417] = 32'b0101000001110000_1_xx_111_xxx_000_0_1_01;
      patterns[418] = 32'b0100000001110000_0_xx_111_000_xxx_1_x_xx;
      patterns[419] = 32'b0000000000000010_1_xx_xxx_xxx_000_0_x_10;
      patterns[420] = 32'b1000000001110100_1_00_111_100_000_0_x_00;
      patterns[421] = 32'b1001000001110100_1_01_111_100_000_0_x_00;
      patterns[422] = 32'b1010000001110100_1_10_111_100_000_0_x_00;
      patterns[423] = 32'b1011000001110100_1_11_111_100_000_0_x_00;
      patterns[424] = 32'b0101000001110000_1_xx_111_xxx_000_0_1_01;
      patterns[425] = 32'b0100000001110000_0_xx_111_000_xxx_1_x_xx;
      patterns[426] = 32'b0000000000000000_1_xx_xxx_xxx_000_0_x_10;
      patterns[427] = 32'b1000000001110101_1_00_111_101_000_0_x_00;
      patterns[428] = 32'b1001000001110101_1_01_111_101_000_0_x_00;
      patterns[429] = 32'b1010000001110101_1_10_111_101_000_0_x_00;
      patterns[430] = 32'b1011000001110101_1_11_111_101_000_0_x_00;
      patterns[431] = 32'b0101000001110000_1_xx_111_xxx_000_0_1_01;
      patterns[432] = 32'b0100000001110000_0_xx_111_000_xxx_1_x_xx;
      patterns[433] = 32'b0000000001100001_1_xx_xxx_xxx_000_0_x_10;
      patterns[434] = 32'b1000000001110110_1_00_111_110_000_0_x_00;
      patterns[435] = 32'b1001000001110110_1_01_111_110_000_0_x_00;
      patterns[436] = 32'b1010000001110110_1_10_111_110_000_0_x_00;
      patterns[437] = 32'b1011000001110110_1_11_111_110_000_0_x_00;
      patterns[438] = 32'b0101000001110000_1_xx_111_xxx_000_0_1_01;
      patterns[439] = 32'b0100000001110000_0_xx_111_000_xxx_1_x_xx;
      patterns[440] = 32'b0000000000000111_1_xx_xxx_xxx_000_0_x_10;
      patterns[441] = 32'b1000000001110111_1_00_111_111_000_0_x_00;
      patterns[442] = 32'b1001000001110111_1_01_111_111_000_0_x_00;
      patterns[443] = 32'b1010000001110111_1_10_111_111_000_0_x_00;
      patterns[444] = 32'b1011000001110111_1_11_111_111_000_0_x_00;
      patterns[445] = 32'b0101000001110000_1_xx_111_xxx_000_0_1_01;
      patterns[446] = 32'b0100000001110000_0_xx_111_000_xxx_1_x_xx;
      patterns[447] = 32'b0000000010101011_1_xx_xxx_xxx_000_0_x_10;
      patterns[448] = 32'b1000000100000000_1_00_000_000_001_0_x_00;
      patterns[449] = 32'b1001000100000000_1_01_000_000_001_0_x_00;
      patterns[450] = 32'b1010000100000000_1_10_000_000_001_0_x_00;
      patterns[451] = 32'b1011000100000000_1_11_000_000_001_0_x_00;
      patterns[452] = 32'b0101000100000000_1_xx_000_xxx_001_0_1_01;
      patterns[453] = 32'b0100000100000000_0_xx_000_001_xxx_1_x_xx;
      patterns[454] = 32'b0000000110010110_1_xx_xxx_xxx_001_0_x_10;
      patterns[455] = 32'b1000000100000001_1_00_000_001_001_0_x_00;
      patterns[456] = 32'b1001000100000001_1_01_000_001_001_0_x_00;
      patterns[457] = 32'b1010000100000001_1_10_000_001_001_0_x_00;
      patterns[458] = 32'b1011000100000001_1_11_000_001_001_0_x_00;
      patterns[459] = 32'b0101000100000000_1_xx_000_xxx_001_0_1_01;
      patterns[460] = 32'b0100000100000000_0_xx_000_001_xxx_1_x_xx;
      patterns[461] = 32'b0000000100111000_1_xx_xxx_xxx_001_0_x_10;
      patterns[462] = 32'b1000000100000010_1_00_000_010_001_0_x_00;
      patterns[463] = 32'b1001000100000010_1_01_000_010_001_0_x_00;
      patterns[464] = 32'b1010000100000010_1_10_000_010_001_0_x_00;
      patterns[465] = 32'b1011000100000010_1_11_000_010_001_0_x_00;
      patterns[466] = 32'b0101000100000000_1_xx_000_xxx_001_0_1_01;
      patterns[467] = 32'b0100000100000000_0_xx_000_001_xxx_1_x_xx;
      patterns[468] = 32'b0000000101000010_1_xx_xxx_xxx_001_0_x_10;
      patterns[469] = 32'b1000000100000011_1_00_000_011_001_0_x_00;
      patterns[470] = 32'b1001000100000011_1_01_000_011_001_0_x_00;
      patterns[471] = 32'b1010000100000011_1_10_000_011_001_0_x_00;
      patterns[472] = 32'b1011000100000011_1_11_000_011_001_0_x_00;
      patterns[473] = 32'b0101000100000000_1_xx_000_xxx_001_0_1_01;
      patterns[474] = 32'b0100000100000000_0_xx_000_001_xxx_1_x_xx;
      patterns[475] = 32'b0000000100001001_1_xx_xxx_xxx_001_0_x_10;
      patterns[476] = 32'b1000000100000100_1_00_000_100_001_0_x_00;
      patterns[477] = 32'b1001000100000100_1_01_000_100_001_0_x_00;
      patterns[478] = 32'b1010000100000100_1_10_000_100_001_0_x_00;
      patterns[479] = 32'b1011000100000100_1_11_000_100_001_0_x_00;
      patterns[480] = 32'b0101000100000000_1_xx_000_xxx_001_0_1_01;
      patterns[481] = 32'b0100000100000000_0_xx_000_001_xxx_1_x_xx;
      patterns[482] = 32'b0000000101010011_1_xx_xxx_xxx_001_0_x_10;
      patterns[483] = 32'b1000000100000101_1_00_000_101_001_0_x_00;
      patterns[484] = 32'b1001000100000101_1_01_000_101_001_0_x_00;
      patterns[485] = 32'b1010000100000101_1_10_000_101_001_0_x_00;
      patterns[486] = 32'b1011000100000101_1_11_000_101_001_0_x_00;
      patterns[487] = 32'b0101000100000000_1_xx_000_xxx_001_0_1_01;
      patterns[488] = 32'b0100000100000000_0_xx_000_001_xxx_1_x_xx;
      patterns[489] = 32'b0000000110001110_1_xx_xxx_xxx_001_0_x_10;
      patterns[490] = 32'b1000000100000110_1_00_000_110_001_0_x_00;
      patterns[491] = 32'b1001000100000110_1_01_000_110_001_0_x_00;
      patterns[492] = 32'b1010000100000110_1_10_000_110_001_0_x_00;
      patterns[493] = 32'b1011000100000110_1_11_000_110_001_0_x_00;
      patterns[494] = 32'b0101000100000000_1_xx_000_xxx_001_0_1_01;
      patterns[495] = 32'b0100000100000000_0_xx_000_001_xxx_1_x_xx;
      patterns[496] = 32'b0000000101101011_1_xx_xxx_xxx_001_0_x_10;
      patterns[497] = 32'b1000000100000111_1_00_000_111_001_0_x_00;
      patterns[498] = 32'b1001000100000111_1_01_000_111_001_0_x_00;
      patterns[499] = 32'b1010000100000111_1_10_000_111_001_0_x_00;
      patterns[500] = 32'b1011000100000111_1_11_000_111_001_0_x_00;
      patterns[501] = 32'b0101000100000000_1_xx_000_xxx_001_0_1_01;
      patterns[502] = 32'b0100000100000000_0_xx_000_001_xxx_1_x_xx;
      patterns[503] = 32'b0000000100111011_1_xx_xxx_xxx_001_0_x_10;
      patterns[504] = 32'b1000000100010000_1_00_001_000_001_0_x_00;
      patterns[505] = 32'b1001000100010000_1_01_001_000_001_0_x_00;
      patterns[506] = 32'b1010000100010000_1_10_001_000_001_0_x_00;
      patterns[507] = 32'b1011000100010000_1_11_001_000_001_0_x_00;
      patterns[508] = 32'b0101000100010000_1_xx_001_xxx_001_0_1_01;
      patterns[509] = 32'b0100000100010000_0_xx_001_001_xxx_1_x_xx;
      patterns[510] = 32'b0000000111100010_1_xx_xxx_xxx_001_0_x_10;
      patterns[511] = 32'b1000000100010001_1_00_001_001_001_0_x_00;
      patterns[512] = 32'b1001000100010001_1_01_001_001_001_0_x_00;
      patterns[513] = 32'b1010000100010001_1_10_001_001_001_0_x_00;
      patterns[514] = 32'b1011000100010001_1_11_001_001_001_0_x_00;
      patterns[515] = 32'b0101000100010000_1_xx_001_xxx_001_0_1_01;
      patterns[516] = 32'b0100000100010000_0_xx_001_001_xxx_1_x_xx;
      patterns[517] = 32'b0000000110011111_1_xx_xxx_xxx_001_0_x_10;
      patterns[518] = 32'b1000000100010010_1_00_001_010_001_0_x_00;
      patterns[519] = 32'b1001000100010010_1_01_001_010_001_0_x_00;
      patterns[520] = 32'b1010000100010010_1_10_001_010_001_0_x_00;
      patterns[521] = 32'b1011000100010010_1_11_001_010_001_0_x_00;
      patterns[522] = 32'b0101000100010000_1_xx_001_xxx_001_0_1_01;
      patterns[523] = 32'b0100000100010000_0_xx_001_001_xxx_1_x_xx;
      patterns[524] = 32'b0000000100011101_1_xx_xxx_xxx_001_0_x_10;
      patterns[525] = 32'b1000000100010011_1_00_001_011_001_0_x_00;
      patterns[526] = 32'b1001000100010011_1_01_001_011_001_0_x_00;
      patterns[527] = 32'b1010000100010011_1_10_001_011_001_0_x_00;
      patterns[528] = 32'b1011000100010011_1_11_001_011_001_0_x_00;
      patterns[529] = 32'b0101000100010000_1_xx_001_xxx_001_0_1_01;
      patterns[530] = 32'b0100000100010000_0_xx_001_001_xxx_1_x_xx;
      patterns[531] = 32'b0000000110101101_1_xx_xxx_xxx_001_0_x_10;
      patterns[532] = 32'b1000000100010100_1_00_001_100_001_0_x_00;
      patterns[533] = 32'b1001000100010100_1_01_001_100_001_0_x_00;
      patterns[534] = 32'b1010000100010100_1_10_001_100_001_0_x_00;
      patterns[535] = 32'b1011000100010100_1_11_001_100_001_0_x_00;
      patterns[536] = 32'b0101000100010000_1_xx_001_xxx_001_0_1_01;
      patterns[537] = 32'b0100000100010000_0_xx_001_001_xxx_1_x_xx;
      patterns[538] = 32'b0000000101110011_1_xx_xxx_xxx_001_0_x_10;
      patterns[539] = 32'b1000000100010101_1_00_001_101_001_0_x_00;
      patterns[540] = 32'b1001000100010101_1_01_001_101_001_0_x_00;
      patterns[541] = 32'b1010000100010101_1_10_001_101_001_0_x_00;
      patterns[542] = 32'b1011000100010101_1_11_001_101_001_0_x_00;
      patterns[543] = 32'b0101000100010000_1_xx_001_xxx_001_0_1_01;
      patterns[544] = 32'b0100000100010000_0_xx_001_001_xxx_1_x_xx;
      patterns[545] = 32'b0000000111110000_1_xx_xxx_xxx_001_0_x_10;
      patterns[546] = 32'b1000000100010110_1_00_001_110_001_0_x_00;
      patterns[547] = 32'b1001000100010110_1_01_001_110_001_0_x_00;
      patterns[548] = 32'b1010000100010110_1_10_001_110_001_0_x_00;
      patterns[549] = 32'b1011000100010110_1_11_001_110_001_0_x_00;
      patterns[550] = 32'b0101000100010000_1_xx_001_xxx_001_0_1_01;
      patterns[551] = 32'b0100000100010000_0_xx_001_001_xxx_1_x_xx;
      patterns[552] = 32'b0000000111110001_1_xx_xxx_xxx_001_0_x_10;
      patterns[553] = 32'b1000000100010111_1_00_001_111_001_0_x_00;
      patterns[554] = 32'b1001000100010111_1_01_001_111_001_0_x_00;
      patterns[555] = 32'b1010000100010111_1_10_001_111_001_0_x_00;
      patterns[556] = 32'b1011000100010111_1_11_001_111_001_0_x_00;
      patterns[557] = 32'b0101000100010000_1_xx_001_xxx_001_0_1_01;
      patterns[558] = 32'b0100000100010000_0_xx_001_001_xxx_1_x_xx;
      patterns[559] = 32'b0000000100001001_1_xx_xxx_xxx_001_0_x_10;
      patterns[560] = 32'b1000000100100000_1_00_010_000_001_0_x_00;
      patterns[561] = 32'b1001000100100000_1_01_010_000_001_0_x_00;
      patterns[562] = 32'b1010000100100000_1_10_010_000_001_0_x_00;
      patterns[563] = 32'b1011000100100000_1_11_010_000_001_0_x_00;
      patterns[564] = 32'b0101000100100000_1_xx_010_xxx_001_0_1_01;
      patterns[565] = 32'b0100000100100000_0_xx_010_001_xxx_1_x_xx;
      patterns[566] = 32'b0000000100001110_1_xx_xxx_xxx_001_0_x_10;
      patterns[567] = 32'b1000000100100001_1_00_010_001_001_0_x_00;
      patterns[568] = 32'b1001000100100001_1_01_010_001_001_0_x_00;
      patterns[569] = 32'b1010000100100001_1_10_010_001_001_0_x_00;
      patterns[570] = 32'b1011000100100001_1_11_010_001_001_0_x_00;
      patterns[571] = 32'b0101000100100000_1_xx_010_xxx_001_0_1_01;
      patterns[572] = 32'b0100000100100000_0_xx_010_001_xxx_1_x_xx;
      patterns[573] = 32'b0000000101011111_1_xx_xxx_xxx_001_0_x_10;
      patterns[574] = 32'b1000000100100010_1_00_010_010_001_0_x_00;
      patterns[575] = 32'b1001000100100010_1_01_010_010_001_0_x_00;
      patterns[576] = 32'b1010000100100010_1_10_010_010_001_0_x_00;
      patterns[577] = 32'b1011000100100010_1_11_010_010_001_0_x_00;
      patterns[578] = 32'b0101000100100000_1_xx_010_xxx_001_0_1_01;
      patterns[579] = 32'b0100000100100000_0_xx_010_001_xxx_1_x_xx;
      patterns[580] = 32'b0000000100011111_1_xx_xxx_xxx_001_0_x_10;
      patterns[581] = 32'b1000000100100011_1_00_010_011_001_0_x_00;
      patterns[582] = 32'b1001000100100011_1_01_010_011_001_0_x_00;
      patterns[583] = 32'b1010000100100011_1_10_010_011_001_0_x_00;
      patterns[584] = 32'b1011000100100011_1_11_010_011_001_0_x_00;
      patterns[585] = 32'b0101000100100000_1_xx_010_xxx_001_0_1_01;
      patterns[586] = 32'b0100000100100000_0_xx_010_001_xxx_1_x_xx;
      patterns[587] = 32'b0000000110010001_1_xx_xxx_xxx_001_0_x_10;
      patterns[588] = 32'b1000000100100100_1_00_010_100_001_0_x_00;
      patterns[589] = 32'b1001000100100100_1_01_010_100_001_0_x_00;
      patterns[590] = 32'b1010000100100100_1_10_010_100_001_0_x_00;
      patterns[591] = 32'b1011000100100100_1_11_010_100_001_0_x_00;
      patterns[592] = 32'b0101000100100000_1_xx_010_xxx_001_0_1_01;
      patterns[593] = 32'b0100000100100000_0_xx_010_001_xxx_1_x_xx;
      patterns[594] = 32'b0000000111111101_1_xx_xxx_xxx_001_0_x_10;
      patterns[595] = 32'b1000000100100101_1_00_010_101_001_0_x_00;
      patterns[596] = 32'b1001000100100101_1_01_010_101_001_0_x_00;
      patterns[597] = 32'b1010000100100101_1_10_010_101_001_0_x_00;
      patterns[598] = 32'b1011000100100101_1_11_010_101_001_0_x_00;
      patterns[599] = 32'b0101000100100000_1_xx_010_xxx_001_0_1_01;
      patterns[600] = 32'b0100000100100000_0_xx_010_001_xxx_1_x_xx;
      patterns[601] = 32'b0000000110101110_1_xx_xxx_xxx_001_0_x_10;
      patterns[602] = 32'b1000000100100110_1_00_010_110_001_0_x_00;
      patterns[603] = 32'b1001000100100110_1_01_010_110_001_0_x_00;
      patterns[604] = 32'b1010000100100110_1_10_010_110_001_0_x_00;
      patterns[605] = 32'b1011000100100110_1_11_010_110_001_0_x_00;
      patterns[606] = 32'b0101000100100000_1_xx_010_xxx_001_0_1_01;
      patterns[607] = 32'b0100000100100000_0_xx_010_001_xxx_1_x_xx;
      patterns[608] = 32'b0000000110001100_1_xx_xxx_xxx_001_0_x_10;
      patterns[609] = 32'b1000000100100111_1_00_010_111_001_0_x_00;
      patterns[610] = 32'b1001000100100111_1_01_010_111_001_0_x_00;
      patterns[611] = 32'b1010000100100111_1_10_010_111_001_0_x_00;
      patterns[612] = 32'b1011000100100111_1_11_010_111_001_0_x_00;
      patterns[613] = 32'b0101000100100000_1_xx_010_xxx_001_0_1_01;
      patterns[614] = 32'b0100000100100000_0_xx_010_001_xxx_1_x_xx;
      patterns[615] = 32'b0000000110111010_1_xx_xxx_xxx_001_0_x_10;
      patterns[616] = 32'b1000000100110000_1_00_011_000_001_0_x_00;
      patterns[617] = 32'b1001000100110000_1_01_011_000_001_0_x_00;
      patterns[618] = 32'b1010000100110000_1_10_011_000_001_0_x_00;
      patterns[619] = 32'b1011000100110000_1_11_011_000_001_0_x_00;
      patterns[620] = 32'b0101000100110000_1_xx_011_xxx_001_0_1_01;
      patterns[621] = 32'b0100000100110000_0_xx_011_001_xxx_1_x_xx;
      patterns[622] = 32'b0000000100001100_1_xx_xxx_xxx_001_0_x_10;
      patterns[623] = 32'b1000000100110001_1_00_011_001_001_0_x_00;
      patterns[624] = 32'b1001000100110001_1_01_011_001_001_0_x_00;
      patterns[625] = 32'b1010000100110001_1_10_011_001_001_0_x_00;
      patterns[626] = 32'b1011000100110001_1_11_011_001_001_0_x_00;
      patterns[627] = 32'b0101000100110000_1_xx_011_xxx_001_0_1_01;
      patterns[628] = 32'b0100000100110000_0_xx_011_001_xxx_1_x_xx;
      patterns[629] = 32'b0000000110000011_1_xx_xxx_xxx_001_0_x_10;
      patterns[630] = 32'b1000000100110010_1_00_011_010_001_0_x_00;
      patterns[631] = 32'b1001000100110010_1_01_011_010_001_0_x_00;
      patterns[632] = 32'b1010000100110010_1_10_011_010_001_0_x_00;
      patterns[633] = 32'b1011000100110010_1_11_011_010_001_0_x_00;
      patterns[634] = 32'b0101000100110000_1_xx_011_xxx_001_0_1_01;
      patterns[635] = 32'b0100000100110000_0_xx_011_001_xxx_1_x_xx;
      patterns[636] = 32'b0000000110110010_1_xx_xxx_xxx_001_0_x_10;
      patterns[637] = 32'b1000000100110011_1_00_011_011_001_0_x_00;
      patterns[638] = 32'b1001000100110011_1_01_011_011_001_0_x_00;
      patterns[639] = 32'b1010000100110011_1_10_011_011_001_0_x_00;
      patterns[640] = 32'b1011000100110011_1_11_011_011_001_0_x_00;
      patterns[641] = 32'b0101000100110000_1_xx_011_xxx_001_0_1_01;
      patterns[642] = 32'b0100000100110000_0_xx_011_001_xxx_1_x_xx;
      patterns[643] = 32'b0000000110110000_1_xx_xxx_xxx_001_0_x_10;
      patterns[644] = 32'b1000000100110100_1_00_011_100_001_0_x_00;
      patterns[645] = 32'b1001000100110100_1_01_011_100_001_0_x_00;
      patterns[646] = 32'b1010000100110100_1_10_011_100_001_0_x_00;
      patterns[647] = 32'b1011000100110100_1_11_011_100_001_0_x_00;
      patterns[648] = 32'b0101000100110000_1_xx_011_xxx_001_0_1_01;
      patterns[649] = 32'b0100000100110000_0_xx_011_001_xxx_1_x_xx;
      patterns[650] = 32'b0000000111101110_1_xx_xxx_xxx_001_0_x_10;
      patterns[651] = 32'b1000000100110101_1_00_011_101_001_0_x_00;
      patterns[652] = 32'b1001000100110101_1_01_011_101_001_0_x_00;
      patterns[653] = 32'b1010000100110101_1_10_011_101_001_0_x_00;
      patterns[654] = 32'b1011000100110101_1_11_011_101_001_0_x_00;
      patterns[655] = 32'b0101000100110000_1_xx_011_xxx_001_0_1_01;
      patterns[656] = 32'b0100000100110000_0_xx_011_001_xxx_1_x_xx;
      patterns[657] = 32'b0000000100111101_1_xx_xxx_xxx_001_0_x_10;
      patterns[658] = 32'b1000000100110110_1_00_011_110_001_0_x_00;
      patterns[659] = 32'b1001000100110110_1_01_011_110_001_0_x_00;
      patterns[660] = 32'b1010000100110110_1_10_011_110_001_0_x_00;
      patterns[661] = 32'b1011000100110110_1_11_011_110_001_0_x_00;
      patterns[662] = 32'b0101000100110000_1_xx_011_xxx_001_0_1_01;
      patterns[663] = 32'b0100000100110000_0_xx_011_001_xxx_1_x_xx;
      patterns[664] = 32'b0000000110001010_1_xx_xxx_xxx_001_0_x_10;
      patterns[665] = 32'b1000000100110111_1_00_011_111_001_0_x_00;
      patterns[666] = 32'b1001000100110111_1_01_011_111_001_0_x_00;
      patterns[667] = 32'b1010000100110111_1_10_011_111_001_0_x_00;
      patterns[668] = 32'b1011000100110111_1_11_011_111_001_0_x_00;
      patterns[669] = 32'b0101000100110000_1_xx_011_xxx_001_0_1_01;
      patterns[670] = 32'b0100000100110000_0_xx_011_001_xxx_1_x_xx;
      patterns[671] = 32'b0000000111001110_1_xx_xxx_xxx_001_0_x_10;
      patterns[672] = 32'b1000000101000000_1_00_100_000_001_0_x_00;
      patterns[673] = 32'b1001000101000000_1_01_100_000_001_0_x_00;
      patterns[674] = 32'b1010000101000000_1_10_100_000_001_0_x_00;
      patterns[675] = 32'b1011000101000000_1_11_100_000_001_0_x_00;
      patterns[676] = 32'b0101000101000000_1_xx_100_xxx_001_0_1_01;
      patterns[677] = 32'b0100000101000000_0_xx_100_001_xxx_1_x_xx;
      patterns[678] = 32'b0000000111111001_1_xx_xxx_xxx_001_0_x_10;
      patterns[679] = 32'b1000000101000001_1_00_100_001_001_0_x_00;
      patterns[680] = 32'b1001000101000001_1_01_100_001_001_0_x_00;
      patterns[681] = 32'b1010000101000001_1_10_100_001_001_0_x_00;
      patterns[682] = 32'b1011000101000001_1_11_100_001_001_0_x_00;
      patterns[683] = 32'b0101000101000000_1_xx_100_xxx_001_0_1_01;
      patterns[684] = 32'b0100000101000000_0_xx_100_001_xxx_1_x_xx;
      patterns[685] = 32'b0000000111110101_1_xx_xxx_xxx_001_0_x_10;
      patterns[686] = 32'b1000000101000010_1_00_100_010_001_0_x_00;
      patterns[687] = 32'b1001000101000010_1_01_100_010_001_0_x_00;
      patterns[688] = 32'b1010000101000010_1_10_100_010_001_0_x_00;
      patterns[689] = 32'b1011000101000010_1_11_100_010_001_0_x_00;
      patterns[690] = 32'b0101000101000000_1_xx_100_xxx_001_0_1_01;
      patterns[691] = 32'b0100000101000000_0_xx_100_001_xxx_1_x_xx;
      patterns[692] = 32'b0000000110011001_1_xx_xxx_xxx_001_0_x_10;
      patterns[693] = 32'b1000000101000011_1_00_100_011_001_0_x_00;
      patterns[694] = 32'b1001000101000011_1_01_100_011_001_0_x_00;
      patterns[695] = 32'b1010000101000011_1_10_100_011_001_0_x_00;
      patterns[696] = 32'b1011000101000011_1_11_100_011_001_0_x_00;
      patterns[697] = 32'b0101000101000000_1_xx_100_xxx_001_0_1_01;
      patterns[698] = 32'b0100000101000000_0_xx_100_001_xxx_1_x_xx;
      patterns[699] = 32'b0000000110100111_1_xx_xxx_xxx_001_0_x_10;
      patterns[700] = 32'b1000000101000100_1_00_100_100_001_0_x_00;
      patterns[701] = 32'b1001000101000100_1_01_100_100_001_0_x_00;
      patterns[702] = 32'b1010000101000100_1_10_100_100_001_0_x_00;
      patterns[703] = 32'b1011000101000100_1_11_100_100_001_0_x_00;
      patterns[704] = 32'b0101000101000000_1_xx_100_xxx_001_0_1_01;
      patterns[705] = 32'b0100000101000000_0_xx_100_001_xxx_1_x_xx;
      patterns[706] = 32'b0000000100111001_1_xx_xxx_xxx_001_0_x_10;
      patterns[707] = 32'b1000000101000101_1_00_100_101_001_0_x_00;
      patterns[708] = 32'b1001000101000101_1_01_100_101_001_0_x_00;
      patterns[709] = 32'b1010000101000101_1_10_100_101_001_0_x_00;
      patterns[710] = 32'b1011000101000101_1_11_100_101_001_0_x_00;
      patterns[711] = 32'b0101000101000000_1_xx_100_xxx_001_0_1_01;
      patterns[712] = 32'b0100000101000000_0_xx_100_001_xxx_1_x_xx;
      patterns[713] = 32'b0000000100101111_1_xx_xxx_xxx_001_0_x_10;
      patterns[714] = 32'b1000000101000110_1_00_100_110_001_0_x_00;
      patterns[715] = 32'b1001000101000110_1_01_100_110_001_0_x_00;
      patterns[716] = 32'b1010000101000110_1_10_100_110_001_0_x_00;
      patterns[717] = 32'b1011000101000110_1_11_100_110_001_0_x_00;
      patterns[718] = 32'b0101000101000000_1_xx_100_xxx_001_0_1_01;
      patterns[719] = 32'b0100000101000000_0_xx_100_001_xxx_1_x_xx;
      patterns[720] = 32'b0000000101110100_1_xx_xxx_xxx_001_0_x_10;
      patterns[721] = 32'b1000000101000111_1_00_100_111_001_0_x_00;
      patterns[722] = 32'b1001000101000111_1_01_100_111_001_0_x_00;
      patterns[723] = 32'b1010000101000111_1_10_100_111_001_0_x_00;
      patterns[724] = 32'b1011000101000111_1_11_100_111_001_0_x_00;
      patterns[725] = 32'b0101000101000000_1_xx_100_xxx_001_0_1_01;
      patterns[726] = 32'b0100000101000000_0_xx_100_001_xxx_1_x_xx;
      patterns[727] = 32'b0000000101111001_1_xx_xxx_xxx_001_0_x_10;
      patterns[728] = 32'b1000000101010000_1_00_101_000_001_0_x_00;
      patterns[729] = 32'b1001000101010000_1_01_101_000_001_0_x_00;
      patterns[730] = 32'b1010000101010000_1_10_101_000_001_0_x_00;
      patterns[731] = 32'b1011000101010000_1_11_101_000_001_0_x_00;
      patterns[732] = 32'b0101000101010000_1_xx_101_xxx_001_0_1_01;
      patterns[733] = 32'b0100000101010000_0_xx_101_001_xxx_1_x_xx;
      patterns[734] = 32'b0000000100110001_1_xx_xxx_xxx_001_0_x_10;
      patterns[735] = 32'b1000000101010001_1_00_101_001_001_0_x_00;
      patterns[736] = 32'b1001000101010001_1_01_101_001_001_0_x_00;
      patterns[737] = 32'b1010000101010001_1_10_101_001_001_0_x_00;
      patterns[738] = 32'b1011000101010001_1_11_101_001_001_0_x_00;
      patterns[739] = 32'b0101000101010000_1_xx_101_xxx_001_0_1_01;
      patterns[740] = 32'b0100000101010000_0_xx_101_001_xxx_1_x_xx;
      patterns[741] = 32'b0000000101110001_1_xx_xxx_xxx_001_0_x_10;
      patterns[742] = 32'b1000000101010010_1_00_101_010_001_0_x_00;
      patterns[743] = 32'b1001000101010010_1_01_101_010_001_0_x_00;
      patterns[744] = 32'b1010000101010010_1_10_101_010_001_0_x_00;
      patterns[745] = 32'b1011000101010010_1_11_101_010_001_0_x_00;
      patterns[746] = 32'b0101000101010000_1_xx_101_xxx_001_0_1_01;
      patterns[747] = 32'b0100000101010000_0_xx_101_001_xxx_1_x_xx;
      patterns[748] = 32'b0000000101100111_1_xx_xxx_xxx_001_0_x_10;
      patterns[749] = 32'b1000000101010011_1_00_101_011_001_0_x_00;
      patterns[750] = 32'b1001000101010011_1_01_101_011_001_0_x_00;
      patterns[751] = 32'b1010000101010011_1_10_101_011_001_0_x_00;
      patterns[752] = 32'b1011000101010011_1_11_101_011_001_0_x_00;
      patterns[753] = 32'b0101000101010000_1_xx_101_xxx_001_0_1_01;
      patterns[754] = 32'b0100000101010000_0_xx_101_001_xxx_1_x_xx;
      patterns[755] = 32'b0000000100111110_1_xx_xxx_xxx_001_0_x_10;
      patterns[756] = 32'b1000000101010100_1_00_101_100_001_0_x_00;
      patterns[757] = 32'b1001000101010100_1_01_101_100_001_0_x_00;
      patterns[758] = 32'b1010000101010100_1_10_101_100_001_0_x_00;
      patterns[759] = 32'b1011000101010100_1_11_101_100_001_0_x_00;
      patterns[760] = 32'b0101000101010000_1_xx_101_xxx_001_0_1_01;
      patterns[761] = 32'b0100000101010000_0_xx_101_001_xxx_1_x_xx;
      patterns[762] = 32'b0000000110011100_1_xx_xxx_xxx_001_0_x_10;
      patterns[763] = 32'b1000000101010101_1_00_101_101_001_0_x_00;
      patterns[764] = 32'b1001000101010101_1_01_101_101_001_0_x_00;
      patterns[765] = 32'b1010000101010101_1_10_101_101_001_0_x_00;
      patterns[766] = 32'b1011000101010101_1_11_101_101_001_0_x_00;
      patterns[767] = 32'b0101000101010000_1_xx_101_xxx_001_0_1_01;
      patterns[768] = 32'b0100000101010000_0_xx_101_001_xxx_1_x_xx;
      patterns[769] = 32'b0000000100011101_1_xx_xxx_xxx_001_0_x_10;
      patterns[770] = 32'b1000000101010110_1_00_101_110_001_0_x_00;
      patterns[771] = 32'b1001000101010110_1_01_101_110_001_0_x_00;
      patterns[772] = 32'b1010000101010110_1_10_101_110_001_0_x_00;
      patterns[773] = 32'b1011000101010110_1_11_101_110_001_0_x_00;
      patterns[774] = 32'b0101000101010000_1_xx_101_xxx_001_0_1_01;
      patterns[775] = 32'b0100000101010000_0_xx_101_001_xxx_1_x_xx;
      patterns[776] = 32'b0000000100111110_1_xx_xxx_xxx_001_0_x_10;
      patterns[777] = 32'b1000000101010111_1_00_101_111_001_0_x_00;
      patterns[778] = 32'b1001000101010111_1_01_101_111_001_0_x_00;
      patterns[779] = 32'b1010000101010111_1_10_101_111_001_0_x_00;
      patterns[780] = 32'b1011000101010111_1_11_101_111_001_0_x_00;
      patterns[781] = 32'b0101000101010000_1_xx_101_xxx_001_0_1_01;
      patterns[782] = 32'b0100000101010000_0_xx_101_001_xxx_1_x_xx;
      patterns[783] = 32'b0000000110100100_1_xx_xxx_xxx_001_0_x_10;
      patterns[784] = 32'b1000000101100000_1_00_110_000_001_0_x_00;
      patterns[785] = 32'b1001000101100000_1_01_110_000_001_0_x_00;
      patterns[786] = 32'b1010000101100000_1_10_110_000_001_0_x_00;
      patterns[787] = 32'b1011000101100000_1_11_110_000_001_0_x_00;
      patterns[788] = 32'b0101000101100000_1_xx_110_xxx_001_0_1_01;
      patterns[789] = 32'b0100000101100000_0_xx_110_001_xxx_1_x_xx;
      patterns[790] = 32'b0000000100101100_1_xx_xxx_xxx_001_0_x_10;
      patterns[791] = 32'b1000000101100001_1_00_110_001_001_0_x_00;
      patterns[792] = 32'b1001000101100001_1_01_110_001_001_0_x_00;
      patterns[793] = 32'b1010000101100001_1_10_110_001_001_0_x_00;
      patterns[794] = 32'b1011000101100001_1_11_110_001_001_0_x_00;
      patterns[795] = 32'b0101000101100000_1_xx_110_xxx_001_0_1_01;
      patterns[796] = 32'b0100000101100000_0_xx_110_001_xxx_1_x_xx;
      patterns[797] = 32'b0000000101001110_1_xx_xxx_xxx_001_0_x_10;
      patterns[798] = 32'b1000000101100010_1_00_110_010_001_0_x_00;
      patterns[799] = 32'b1001000101100010_1_01_110_010_001_0_x_00;
      patterns[800] = 32'b1010000101100010_1_10_110_010_001_0_x_00;
      patterns[801] = 32'b1011000101100010_1_11_110_010_001_0_x_00;
      patterns[802] = 32'b0101000101100000_1_xx_110_xxx_001_0_1_01;
      patterns[803] = 32'b0100000101100000_0_xx_110_001_xxx_1_x_xx;
      patterns[804] = 32'b0000000100000001_1_xx_xxx_xxx_001_0_x_10;
      patterns[805] = 32'b1000000101100011_1_00_110_011_001_0_x_00;
      patterns[806] = 32'b1001000101100011_1_01_110_011_001_0_x_00;
      patterns[807] = 32'b1010000101100011_1_10_110_011_001_0_x_00;
      patterns[808] = 32'b1011000101100011_1_11_110_011_001_0_x_00;
      patterns[809] = 32'b0101000101100000_1_xx_110_xxx_001_0_1_01;
      patterns[810] = 32'b0100000101100000_0_xx_110_001_xxx_1_x_xx;
      patterns[811] = 32'b0000000101010000_1_xx_xxx_xxx_001_0_x_10;
      patterns[812] = 32'b1000000101100100_1_00_110_100_001_0_x_00;
      patterns[813] = 32'b1001000101100100_1_01_110_100_001_0_x_00;
      patterns[814] = 32'b1010000101100100_1_10_110_100_001_0_x_00;
      patterns[815] = 32'b1011000101100100_1_11_110_100_001_0_x_00;
      patterns[816] = 32'b0101000101100000_1_xx_110_xxx_001_0_1_01;
      patterns[817] = 32'b0100000101100000_0_xx_110_001_xxx_1_x_xx;
      patterns[818] = 32'b0000000110101000_1_xx_xxx_xxx_001_0_x_10;
      patterns[819] = 32'b1000000101100101_1_00_110_101_001_0_x_00;
      patterns[820] = 32'b1001000101100101_1_01_110_101_001_0_x_00;
      patterns[821] = 32'b1010000101100101_1_10_110_101_001_0_x_00;
      patterns[822] = 32'b1011000101100101_1_11_110_101_001_0_x_00;
      patterns[823] = 32'b0101000101100000_1_xx_110_xxx_001_0_1_01;
      patterns[824] = 32'b0100000101100000_0_xx_110_001_xxx_1_x_xx;
      patterns[825] = 32'b0000000101110101_1_xx_xxx_xxx_001_0_x_10;
      patterns[826] = 32'b1000000101100110_1_00_110_110_001_0_x_00;
      patterns[827] = 32'b1001000101100110_1_01_110_110_001_0_x_00;
      patterns[828] = 32'b1010000101100110_1_10_110_110_001_0_x_00;
      patterns[829] = 32'b1011000101100110_1_11_110_110_001_0_x_00;
      patterns[830] = 32'b0101000101100000_1_xx_110_xxx_001_0_1_01;
      patterns[831] = 32'b0100000101100000_0_xx_110_001_xxx_1_x_xx;
      patterns[832] = 32'b0000000100001001_1_xx_xxx_xxx_001_0_x_10;
      patterns[833] = 32'b1000000101100111_1_00_110_111_001_0_x_00;
      patterns[834] = 32'b1001000101100111_1_01_110_111_001_0_x_00;
      patterns[835] = 32'b1010000101100111_1_10_110_111_001_0_x_00;
      patterns[836] = 32'b1011000101100111_1_11_110_111_001_0_x_00;
      patterns[837] = 32'b0101000101100000_1_xx_110_xxx_001_0_1_01;
      patterns[838] = 32'b0100000101100000_0_xx_110_001_xxx_1_x_xx;
      patterns[839] = 32'b0000000111010001_1_xx_xxx_xxx_001_0_x_10;
      patterns[840] = 32'b1000000101110000_1_00_111_000_001_0_x_00;
      patterns[841] = 32'b1001000101110000_1_01_111_000_001_0_x_00;
      patterns[842] = 32'b1010000101110000_1_10_111_000_001_0_x_00;
      patterns[843] = 32'b1011000101110000_1_11_111_000_001_0_x_00;
      patterns[844] = 32'b0101000101110000_1_xx_111_xxx_001_0_1_01;
      patterns[845] = 32'b0100000101110000_0_xx_111_001_xxx_1_x_xx;
      patterns[846] = 32'b0000000110101111_1_xx_xxx_xxx_001_0_x_10;
      patterns[847] = 32'b1000000101110001_1_00_111_001_001_0_x_00;
      patterns[848] = 32'b1001000101110001_1_01_111_001_001_0_x_00;
      patterns[849] = 32'b1010000101110001_1_10_111_001_001_0_x_00;
      patterns[850] = 32'b1011000101110001_1_11_111_001_001_0_x_00;
      patterns[851] = 32'b0101000101110000_1_xx_111_xxx_001_0_1_01;
      patterns[852] = 32'b0100000101110000_0_xx_111_001_xxx_1_x_xx;
      patterns[853] = 32'b0000000110101101_1_xx_xxx_xxx_001_0_x_10;
      patterns[854] = 32'b1000000101110010_1_00_111_010_001_0_x_00;
      patterns[855] = 32'b1001000101110010_1_01_111_010_001_0_x_00;
      patterns[856] = 32'b1010000101110010_1_10_111_010_001_0_x_00;
      patterns[857] = 32'b1011000101110010_1_11_111_010_001_0_x_00;
      patterns[858] = 32'b0101000101110000_1_xx_111_xxx_001_0_1_01;
      patterns[859] = 32'b0100000101110000_0_xx_111_001_xxx_1_x_xx;
      patterns[860] = 32'b0000000111110001_1_xx_xxx_xxx_001_0_x_10;
      patterns[861] = 32'b1000000101110011_1_00_111_011_001_0_x_00;
      patterns[862] = 32'b1001000101110011_1_01_111_011_001_0_x_00;
      patterns[863] = 32'b1010000101110011_1_10_111_011_001_0_x_00;
      patterns[864] = 32'b1011000101110011_1_11_111_011_001_0_x_00;
      patterns[865] = 32'b0101000101110000_1_xx_111_xxx_001_0_1_01;
      patterns[866] = 32'b0100000101110000_0_xx_111_001_xxx_1_x_xx;
      patterns[867] = 32'b0000000101101111_1_xx_xxx_xxx_001_0_x_10;
      patterns[868] = 32'b1000000101110100_1_00_111_100_001_0_x_00;
      patterns[869] = 32'b1001000101110100_1_01_111_100_001_0_x_00;
      patterns[870] = 32'b1010000101110100_1_10_111_100_001_0_x_00;
      patterns[871] = 32'b1011000101110100_1_11_111_100_001_0_x_00;
      patterns[872] = 32'b0101000101110000_1_xx_111_xxx_001_0_1_01;
      patterns[873] = 32'b0100000101110000_0_xx_111_001_xxx_1_x_xx;
      patterns[874] = 32'b0000000100010110_1_xx_xxx_xxx_001_0_x_10;
      patterns[875] = 32'b1000000101110101_1_00_111_101_001_0_x_00;
      patterns[876] = 32'b1001000101110101_1_01_111_101_001_0_x_00;
      patterns[877] = 32'b1010000101110101_1_10_111_101_001_0_x_00;
      patterns[878] = 32'b1011000101110101_1_11_111_101_001_0_x_00;
      patterns[879] = 32'b0101000101110000_1_xx_111_xxx_001_0_1_01;
      patterns[880] = 32'b0100000101110000_0_xx_111_001_xxx_1_x_xx;
      patterns[881] = 32'b0000000101111110_1_xx_xxx_xxx_001_0_x_10;
      patterns[882] = 32'b1000000101110110_1_00_111_110_001_0_x_00;
      patterns[883] = 32'b1001000101110110_1_01_111_110_001_0_x_00;
      patterns[884] = 32'b1010000101110110_1_10_111_110_001_0_x_00;
      patterns[885] = 32'b1011000101110110_1_11_111_110_001_0_x_00;
      patterns[886] = 32'b0101000101110000_1_xx_111_xxx_001_0_1_01;
      patterns[887] = 32'b0100000101110000_0_xx_111_001_xxx_1_x_xx;
      patterns[888] = 32'b0000000111010101_1_xx_xxx_xxx_001_0_x_10;
      patterns[889] = 32'b1000000101110111_1_00_111_111_001_0_x_00;
      patterns[890] = 32'b1001000101110111_1_01_111_111_001_0_x_00;
      patterns[891] = 32'b1010000101110111_1_10_111_111_001_0_x_00;
      patterns[892] = 32'b1011000101110111_1_11_111_111_001_0_x_00;
      patterns[893] = 32'b0101000101110000_1_xx_111_xxx_001_0_1_01;
      patterns[894] = 32'b0100000101110000_0_xx_111_001_xxx_1_x_xx;
      patterns[895] = 32'b0000000111101100_1_xx_xxx_xxx_001_0_x_10;
      patterns[896] = 32'b1000001000000000_1_00_000_000_010_0_x_00;
      patterns[897] = 32'b1001001000000000_1_01_000_000_010_0_x_00;
      patterns[898] = 32'b1010001000000000_1_10_000_000_010_0_x_00;
      patterns[899] = 32'b1011001000000000_1_11_000_000_010_0_x_00;
      patterns[900] = 32'b0101001000000000_1_xx_000_xxx_010_0_1_01;
      patterns[901] = 32'b0100001000000000_0_xx_000_010_xxx_1_x_xx;
      patterns[902] = 32'b0000001000100011_1_xx_xxx_xxx_010_0_x_10;
      patterns[903] = 32'b1000001000000001_1_00_000_001_010_0_x_00;
      patterns[904] = 32'b1001001000000001_1_01_000_001_010_0_x_00;
      patterns[905] = 32'b1010001000000001_1_10_000_001_010_0_x_00;
      patterns[906] = 32'b1011001000000001_1_11_000_001_010_0_x_00;
      patterns[907] = 32'b0101001000000000_1_xx_000_xxx_010_0_1_01;
      patterns[908] = 32'b0100001000000000_0_xx_000_010_xxx_1_x_xx;
      patterns[909] = 32'b0000001011100011_1_xx_xxx_xxx_010_0_x_10;
      patterns[910] = 32'b1000001000000010_1_00_000_010_010_0_x_00;
      patterns[911] = 32'b1001001000000010_1_01_000_010_010_0_x_00;
      patterns[912] = 32'b1010001000000010_1_10_000_010_010_0_x_00;
      patterns[913] = 32'b1011001000000010_1_11_000_010_010_0_x_00;
      patterns[914] = 32'b0101001000000000_1_xx_000_xxx_010_0_1_01;
      patterns[915] = 32'b0100001000000000_0_xx_000_010_xxx_1_x_xx;
      patterns[916] = 32'b0000001010110000_1_xx_xxx_xxx_010_0_x_10;
      patterns[917] = 32'b1000001000000011_1_00_000_011_010_0_x_00;
      patterns[918] = 32'b1001001000000011_1_01_000_011_010_0_x_00;
      patterns[919] = 32'b1010001000000011_1_10_000_011_010_0_x_00;
      patterns[920] = 32'b1011001000000011_1_11_000_011_010_0_x_00;
      patterns[921] = 32'b0101001000000000_1_xx_000_xxx_010_0_1_01;
      patterns[922] = 32'b0100001000000000_0_xx_000_010_xxx_1_x_xx;
      patterns[923] = 32'b0000001011100101_1_xx_xxx_xxx_010_0_x_10;
      patterns[924] = 32'b1000001000000100_1_00_000_100_010_0_x_00;
      patterns[925] = 32'b1001001000000100_1_01_000_100_010_0_x_00;
      patterns[926] = 32'b1010001000000100_1_10_000_100_010_0_x_00;
      patterns[927] = 32'b1011001000000100_1_11_000_100_010_0_x_00;
      patterns[928] = 32'b0101001000000000_1_xx_000_xxx_010_0_1_01;
      patterns[929] = 32'b0100001000000000_0_xx_000_010_xxx_1_x_xx;
      patterns[930] = 32'b0000001011010111_1_xx_xxx_xxx_010_0_x_10;
      patterns[931] = 32'b1000001000000101_1_00_000_101_010_0_x_00;
      patterns[932] = 32'b1001001000000101_1_01_000_101_010_0_x_00;
      patterns[933] = 32'b1010001000000101_1_10_000_101_010_0_x_00;
      patterns[934] = 32'b1011001000000101_1_11_000_101_010_0_x_00;
      patterns[935] = 32'b0101001000000000_1_xx_000_xxx_010_0_1_01;
      patterns[936] = 32'b0100001000000000_0_xx_000_010_xxx_1_x_xx;
      patterns[937] = 32'b0000001011100111_1_xx_xxx_xxx_010_0_x_10;
      patterns[938] = 32'b1000001000000110_1_00_000_110_010_0_x_00;
      patterns[939] = 32'b1001001000000110_1_01_000_110_010_0_x_00;
      patterns[940] = 32'b1010001000000110_1_10_000_110_010_0_x_00;
      patterns[941] = 32'b1011001000000110_1_11_000_110_010_0_x_00;
      patterns[942] = 32'b0101001000000000_1_xx_000_xxx_010_0_1_01;
      patterns[943] = 32'b0100001000000000_0_xx_000_010_xxx_1_x_xx;
      patterns[944] = 32'b0000001011110100_1_xx_xxx_xxx_010_0_x_10;
      patterns[945] = 32'b1000001000000111_1_00_000_111_010_0_x_00;
      patterns[946] = 32'b1001001000000111_1_01_000_111_010_0_x_00;
      patterns[947] = 32'b1010001000000111_1_10_000_111_010_0_x_00;
      patterns[948] = 32'b1011001000000111_1_11_000_111_010_0_x_00;
      patterns[949] = 32'b0101001000000000_1_xx_000_xxx_010_0_1_01;
      patterns[950] = 32'b0100001000000000_0_xx_000_010_xxx_1_x_xx;
      patterns[951] = 32'b0000001000101011_1_xx_xxx_xxx_010_0_x_10;
      patterns[952] = 32'b1000001000010000_1_00_001_000_010_0_x_00;
      patterns[953] = 32'b1001001000010000_1_01_001_000_010_0_x_00;
      patterns[954] = 32'b1010001000010000_1_10_001_000_010_0_x_00;
      patterns[955] = 32'b1011001000010000_1_11_001_000_010_0_x_00;
      patterns[956] = 32'b0101001000010000_1_xx_001_xxx_010_0_1_01;
      patterns[957] = 32'b0100001000010000_0_xx_001_010_xxx_1_x_xx;
      patterns[958] = 32'b0000001000001001_1_xx_xxx_xxx_010_0_x_10;
      patterns[959] = 32'b1000001000010001_1_00_001_001_010_0_x_00;
      patterns[960] = 32'b1001001000010001_1_01_001_001_010_0_x_00;
      patterns[961] = 32'b1010001000010001_1_10_001_001_010_0_x_00;
      patterns[962] = 32'b1011001000010001_1_11_001_001_010_0_x_00;
      patterns[963] = 32'b0101001000010000_1_xx_001_xxx_010_0_1_01;
      patterns[964] = 32'b0100001000010000_0_xx_001_010_xxx_1_x_xx;
      patterns[965] = 32'b0000001000011101_1_xx_xxx_xxx_010_0_x_10;
      patterns[966] = 32'b1000001000010010_1_00_001_010_010_0_x_00;
      patterns[967] = 32'b1001001000010010_1_01_001_010_010_0_x_00;
      patterns[968] = 32'b1010001000010010_1_10_001_010_010_0_x_00;
      patterns[969] = 32'b1011001000010010_1_11_001_010_010_0_x_00;
      patterns[970] = 32'b0101001000010000_1_xx_001_xxx_010_0_1_01;
      patterns[971] = 32'b0100001000010000_0_xx_001_010_xxx_1_x_xx;
      patterns[972] = 32'b0000001000110000_1_xx_xxx_xxx_010_0_x_10;
      patterns[973] = 32'b1000001000010011_1_00_001_011_010_0_x_00;
      patterns[974] = 32'b1001001000010011_1_01_001_011_010_0_x_00;
      patterns[975] = 32'b1010001000010011_1_10_001_011_010_0_x_00;
      patterns[976] = 32'b1011001000010011_1_11_001_011_010_0_x_00;
      patterns[977] = 32'b0101001000010000_1_xx_001_xxx_010_0_1_01;
      patterns[978] = 32'b0100001000010000_0_xx_001_010_xxx_1_x_xx;
      patterns[979] = 32'b0000001011100010_1_xx_xxx_xxx_010_0_x_10;
      patterns[980] = 32'b1000001000010100_1_00_001_100_010_0_x_00;
      patterns[981] = 32'b1001001000010100_1_01_001_100_010_0_x_00;
      patterns[982] = 32'b1010001000010100_1_10_001_100_010_0_x_00;
      patterns[983] = 32'b1011001000010100_1_11_001_100_010_0_x_00;
      patterns[984] = 32'b0101001000010000_1_xx_001_xxx_010_0_1_01;
      patterns[985] = 32'b0100001000010000_0_xx_001_010_xxx_1_x_xx;
      patterns[986] = 32'b0000001001111100_1_xx_xxx_xxx_010_0_x_10;
      patterns[987] = 32'b1000001000010101_1_00_001_101_010_0_x_00;
      patterns[988] = 32'b1001001000010101_1_01_001_101_010_0_x_00;
      patterns[989] = 32'b1010001000010101_1_10_001_101_010_0_x_00;
      patterns[990] = 32'b1011001000010101_1_11_001_101_010_0_x_00;
      patterns[991] = 32'b0101001000010000_1_xx_001_xxx_010_0_1_01;
      patterns[992] = 32'b0100001000010000_0_xx_001_010_xxx_1_x_xx;
      patterns[993] = 32'b0000001010010100_1_xx_xxx_xxx_010_0_x_10;
      patterns[994] = 32'b1000001000010110_1_00_001_110_010_0_x_00;
      patterns[995] = 32'b1001001000010110_1_01_001_110_010_0_x_00;
      patterns[996] = 32'b1010001000010110_1_10_001_110_010_0_x_00;
      patterns[997] = 32'b1011001000010110_1_11_001_110_010_0_x_00;
      patterns[998] = 32'b0101001000010000_1_xx_001_xxx_010_0_1_01;
      patterns[999] = 32'b0100001000010000_0_xx_001_010_xxx_1_x_xx;
      patterns[1000] = 32'b0000001000010100_1_xx_xxx_xxx_010_0_x_10;
      patterns[1001] = 32'b1000001000010111_1_00_001_111_010_0_x_00;
      patterns[1002] = 32'b1001001000010111_1_01_001_111_010_0_x_00;
      patterns[1003] = 32'b1010001000010111_1_10_001_111_010_0_x_00;
      patterns[1004] = 32'b1011001000010111_1_11_001_111_010_0_x_00;
      patterns[1005] = 32'b0101001000010000_1_xx_001_xxx_010_0_1_01;
      patterns[1006] = 32'b0100001000010000_0_xx_001_010_xxx_1_x_xx;
      patterns[1007] = 32'b0000001010011010_1_xx_xxx_xxx_010_0_x_10;
      patterns[1008] = 32'b1000001000100000_1_00_010_000_010_0_x_00;
      patterns[1009] = 32'b1001001000100000_1_01_010_000_010_0_x_00;
      patterns[1010] = 32'b1010001000100000_1_10_010_000_010_0_x_00;
      patterns[1011] = 32'b1011001000100000_1_11_010_000_010_0_x_00;
      patterns[1012] = 32'b0101001000100000_1_xx_010_xxx_010_0_1_01;
      patterns[1013] = 32'b0100001000100000_0_xx_010_010_xxx_1_x_xx;
      patterns[1014] = 32'b0000001011001101_1_xx_xxx_xxx_010_0_x_10;
      patterns[1015] = 32'b1000001000100001_1_00_010_001_010_0_x_00;
      patterns[1016] = 32'b1001001000100001_1_01_010_001_010_0_x_00;
      patterns[1017] = 32'b1010001000100001_1_10_010_001_010_0_x_00;
      patterns[1018] = 32'b1011001000100001_1_11_010_001_010_0_x_00;
      patterns[1019] = 32'b0101001000100000_1_xx_010_xxx_010_0_1_01;
      patterns[1020] = 32'b0100001000100000_0_xx_010_010_xxx_1_x_xx;
      patterns[1021] = 32'b0000001010010000_1_xx_xxx_xxx_010_0_x_10;
      patterns[1022] = 32'b1000001000100010_1_00_010_010_010_0_x_00;
      patterns[1023] = 32'b1001001000100010_1_01_010_010_010_0_x_00;
      patterns[1024] = 32'b1010001000100010_1_10_010_010_010_0_x_00;
      patterns[1025] = 32'b1011001000100010_1_11_010_010_010_0_x_00;
      patterns[1026] = 32'b0101001000100000_1_xx_010_xxx_010_0_1_01;
      patterns[1027] = 32'b0100001000100000_0_xx_010_010_xxx_1_x_xx;
      patterns[1028] = 32'b0000001001000100_1_xx_xxx_xxx_010_0_x_10;
      patterns[1029] = 32'b1000001000100011_1_00_010_011_010_0_x_00;
      patterns[1030] = 32'b1001001000100011_1_01_010_011_010_0_x_00;
      patterns[1031] = 32'b1010001000100011_1_10_010_011_010_0_x_00;
      patterns[1032] = 32'b1011001000100011_1_11_010_011_010_0_x_00;
      patterns[1033] = 32'b0101001000100000_1_xx_010_xxx_010_0_1_01;
      patterns[1034] = 32'b0100001000100000_0_xx_010_010_xxx_1_x_xx;
      patterns[1035] = 32'b0000001000000101_1_xx_xxx_xxx_010_0_x_10;
      patterns[1036] = 32'b1000001000100100_1_00_010_100_010_0_x_00;
      patterns[1037] = 32'b1001001000100100_1_01_010_100_010_0_x_00;
      patterns[1038] = 32'b1010001000100100_1_10_010_100_010_0_x_00;
      patterns[1039] = 32'b1011001000100100_1_11_010_100_010_0_x_00;
      patterns[1040] = 32'b0101001000100000_1_xx_010_xxx_010_0_1_01;
      patterns[1041] = 32'b0100001000100000_0_xx_010_010_xxx_1_x_xx;
      patterns[1042] = 32'b0000001011100100_1_xx_xxx_xxx_010_0_x_10;
      patterns[1043] = 32'b1000001000100101_1_00_010_101_010_0_x_00;
      patterns[1044] = 32'b1001001000100101_1_01_010_101_010_0_x_00;
      patterns[1045] = 32'b1010001000100101_1_10_010_101_010_0_x_00;
      patterns[1046] = 32'b1011001000100101_1_11_010_101_010_0_x_00;
      patterns[1047] = 32'b0101001000100000_1_xx_010_xxx_010_0_1_01;
      patterns[1048] = 32'b0100001000100000_0_xx_010_010_xxx_1_x_xx;
      patterns[1049] = 32'b0000001010011000_1_xx_xxx_xxx_010_0_x_10;
      patterns[1050] = 32'b1000001000100110_1_00_010_110_010_0_x_00;
      patterns[1051] = 32'b1001001000100110_1_01_010_110_010_0_x_00;
      patterns[1052] = 32'b1010001000100110_1_10_010_110_010_0_x_00;
      patterns[1053] = 32'b1011001000100110_1_11_010_110_010_0_x_00;
      patterns[1054] = 32'b0101001000100000_1_xx_010_xxx_010_0_1_01;
      patterns[1055] = 32'b0100001000100000_0_xx_010_010_xxx_1_x_xx;
      patterns[1056] = 32'b0000001000110101_1_xx_xxx_xxx_010_0_x_10;
      patterns[1057] = 32'b1000001000100111_1_00_010_111_010_0_x_00;
      patterns[1058] = 32'b1001001000100111_1_01_010_111_010_0_x_00;
      patterns[1059] = 32'b1010001000100111_1_10_010_111_010_0_x_00;
      patterns[1060] = 32'b1011001000100111_1_11_010_111_010_0_x_00;
      patterns[1061] = 32'b0101001000100000_1_xx_010_xxx_010_0_1_01;
      patterns[1062] = 32'b0100001000100000_0_xx_010_010_xxx_1_x_xx;
      patterns[1063] = 32'b0000001011110011_1_xx_xxx_xxx_010_0_x_10;
      patterns[1064] = 32'b1000001000110000_1_00_011_000_010_0_x_00;
      patterns[1065] = 32'b1001001000110000_1_01_011_000_010_0_x_00;
      patterns[1066] = 32'b1010001000110000_1_10_011_000_010_0_x_00;
      patterns[1067] = 32'b1011001000110000_1_11_011_000_010_0_x_00;
      patterns[1068] = 32'b0101001000110000_1_xx_011_xxx_010_0_1_01;
      patterns[1069] = 32'b0100001000110000_0_xx_011_010_xxx_1_x_xx;
      patterns[1070] = 32'b0000001010010111_1_xx_xxx_xxx_010_0_x_10;
      patterns[1071] = 32'b1000001000110001_1_00_011_001_010_0_x_00;
      patterns[1072] = 32'b1001001000110001_1_01_011_001_010_0_x_00;
      patterns[1073] = 32'b1010001000110001_1_10_011_001_010_0_x_00;
      patterns[1074] = 32'b1011001000110001_1_11_011_001_010_0_x_00;
      patterns[1075] = 32'b0101001000110000_1_xx_011_xxx_010_0_1_01;
      patterns[1076] = 32'b0100001000110000_0_xx_011_010_xxx_1_x_xx;
      patterns[1077] = 32'b0000001011001001_1_xx_xxx_xxx_010_0_x_10;
      patterns[1078] = 32'b1000001000110010_1_00_011_010_010_0_x_00;
      patterns[1079] = 32'b1001001000110010_1_01_011_010_010_0_x_00;
      patterns[1080] = 32'b1010001000110010_1_10_011_010_010_0_x_00;
      patterns[1081] = 32'b1011001000110010_1_11_011_010_010_0_x_00;
      patterns[1082] = 32'b0101001000110000_1_xx_011_xxx_010_0_1_01;
      patterns[1083] = 32'b0100001000110000_0_xx_011_010_xxx_1_x_xx;
      patterns[1084] = 32'b0000001010110110_1_xx_xxx_xxx_010_0_x_10;
      patterns[1085] = 32'b1000001000110011_1_00_011_011_010_0_x_00;
      patterns[1086] = 32'b1001001000110011_1_01_011_011_010_0_x_00;
      patterns[1087] = 32'b1010001000110011_1_10_011_011_010_0_x_00;
      patterns[1088] = 32'b1011001000110011_1_11_011_011_010_0_x_00;
      patterns[1089] = 32'b0101001000110000_1_xx_011_xxx_010_0_1_01;
      patterns[1090] = 32'b0100001000110000_0_xx_011_010_xxx_1_x_xx;
      patterns[1091] = 32'b0000001010010010_1_xx_xxx_xxx_010_0_x_10;
      patterns[1092] = 32'b1000001000110100_1_00_011_100_010_0_x_00;
      patterns[1093] = 32'b1001001000110100_1_01_011_100_010_0_x_00;
      patterns[1094] = 32'b1010001000110100_1_10_011_100_010_0_x_00;
      patterns[1095] = 32'b1011001000110100_1_11_011_100_010_0_x_00;
      patterns[1096] = 32'b0101001000110000_1_xx_011_xxx_010_0_1_01;
      patterns[1097] = 32'b0100001000110000_0_xx_011_010_xxx_1_x_xx;
      patterns[1098] = 32'b0000001001001100_1_xx_xxx_xxx_010_0_x_10;
      patterns[1099] = 32'b1000001000110101_1_00_011_101_010_0_x_00;
      patterns[1100] = 32'b1001001000110101_1_01_011_101_010_0_x_00;
      patterns[1101] = 32'b1010001000110101_1_10_011_101_010_0_x_00;
      patterns[1102] = 32'b1011001000110101_1_11_011_101_010_0_x_00;
      patterns[1103] = 32'b0101001000110000_1_xx_011_xxx_010_0_1_01;
      patterns[1104] = 32'b0100001000110000_0_xx_011_010_xxx_1_x_xx;
      patterns[1105] = 32'b0000001010001011_1_xx_xxx_xxx_010_0_x_10;
      patterns[1106] = 32'b1000001000110110_1_00_011_110_010_0_x_00;
      patterns[1107] = 32'b1001001000110110_1_01_011_110_010_0_x_00;
      patterns[1108] = 32'b1010001000110110_1_10_011_110_010_0_x_00;
      patterns[1109] = 32'b1011001000110110_1_11_011_110_010_0_x_00;
      patterns[1110] = 32'b0101001000110000_1_xx_011_xxx_010_0_1_01;
      patterns[1111] = 32'b0100001000110000_0_xx_011_010_xxx_1_x_xx;
      patterns[1112] = 32'b0000001011100111_1_xx_xxx_xxx_010_0_x_10;
      patterns[1113] = 32'b1000001000110111_1_00_011_111_010_0_x_00;
      patterns[1114] = 32'b1001001000110111_1_01_011_111_010_0_x_00;
      patterns[1115] = 32'b1010001000110111_1_10_011_111_010_0_x_00;
      patterns[1116] = 32'b1011001000110111_1_11_011_111_010_0_x_00;
      patterns[1117] = 32'b0101001000110000_1_xx_011_xxx_010_0_1_01;
      patterns[1118] = 32'b0100001000110000_0_xx_011_010_xxx_1_x_xx;
      patterns[1119] = 32'b0000001011010111_1_xx_xxx_xxx_010_0_x_10;
      patterns[1120] = 32'b1000001001000000_1_00_100_000_010_0_x_00;
      patterns[1121] = 32'b1001001001000000_1_01_100_000_010_0_x_00;
      patterns[1122] = 32'b1010001001000000_1_10_100_000_010_0_x_00;
      patterns[1123] = 32'b1011001001000000_1_11_100_000_010_0_x_00;
      patterns[1124] = 32'b0101001001000000_1_xx_100_xxx_010_0_1_01;
      patterns[1125] = 32'b0100001001000000_0_xx_100_010_xxx_1_x_xx;
      patterns[1126] = 32'b0000001010110110_1_xx_xxx_xxx_010_0_x_10;
      patterns[1127] = 32'b1000001001000001_1_00_100_001_010_0_x_00;
      patterns[1128] = 32'b1001001001000001_1_01_100_001_010_0_x_00;
      patterns[1129] = 32'b1010001001000001_1_10_100_001_010_0_x_00;
      patterns[1130] = 32'b1011001001000001_1_11_100_001_010_0_x_00;
      patterns[1131] = 32'b0101001001000000_1_xx_100_xxx_010_0_1_01;
      patterns[1132] = 32'b0100001001000000_0_xx_100_010_xxx_1_x_xx;
      patterns[1133] = 32'b0000001011100011_1_xx_xxx_xxx_010_0_x_10;
      patterns[1134] = 32'b1000001001000010_1_00_100_010_010_0_x_00;
      patterns[1135] = 32'b1001001001000010_1_01_100_010_010_0_x_00;
      patterns[1136] = 32'b1010001001000010_1_10_100_010_010_0_x_00;
      patterns[1137] = 32'b1011001001000010_1_11_100_010_010_0_x_00;
      patterns[1138] = 32'b0101001001000000_1_xx_100_xxx_010_0_1_01;
      patterns[1139] = 32'b0100001001000000_0_xx_100_010_xxx_1_x_xx;
      patterns[1140] = 32'b0000001000011011_1_xx_xxx_xxx_010_0_x_10;
      patterns[1141] = 32'b1000001001000011_1_00_100_011_010_0_x_00;
      patterns[1142] = 32'b1001001001000011_1_01_100_011_010_0_x_00;
      patterns[1143] = 32'b1010001001000011_1_10_100_011_010_0_x_00;
      patterns[1144] = 32'b1011001001000011_1_11_100_011_010_0_x_00;
      patterns[1145] = 32'b0101001001000000_1_xx_100_xxx_010_0_1_01;
      patterns[1146] = 32'b0100001001000000_0_xx_100_010_xxx_1_x_xx;
      patterns[1147] = 32'b0000001011110011_1_xx_xxx_xxx_010_0_x_10;
      patterns[1148] = 32'b1000001001000100_1_00_100_100_010_0_x_00;
      patterns[1149] = 32'b1001001001000100_1_01_100_100_010_0_x_00;
      patterns[1150] = 32'b1010001001000100_1_10_100_100_010_0_x_00;
      patterns[1151] = 32'b1011001001000100_1_11_100_100_010_0_x_00;
      patterns[1152] = 32'b0101001001000000_1_xx_100_xxx_010_0_1_01;
      patterns[1153] = 32'b0100001001000000_0_xx_100_010_xxx_1_x_xx;
      patterns[1154] = 32'b0000001000101011_1_xx_xxx_xxx_010_0_x_10;
      patterns[1155] = 32'b1000001001000101_1_00_100_101_010_0_x_00;
      patterns[1156] = 32'b1001001001000101_1_01_100_101_010_0_x_00;
      patterns[1157] = 32'b1010001001000101_1_10_100_101_010_0_x_00;
      patterns[1158] = 32'b1011001001000101_1_11_100_101_010_0_x_00;
      patterns[1159] = 32'b0101001001000000_1_xx_100_xxx_010_0_1_01;
      patterns[1160] = 32'b0100001001000000_0_xx_100_010_xxx_1_x_xx;
      patterns[1161] = 32'b0000001010100100_1_xx_xxx_xxx_010_0_x_10;
      patterns[1162] = 32'b1000001001000110_1_00_100_110_010_0_x_00;
      patterns[1163] = 32'b1001001001000110_1_01_100_110_010_0_x_00;
      patterns[1164] = 32'b1010001001000110_1_10_100_110_010_0_x_00;
      patterns[1165] = 32'b1011001001000110_1_11_100_110_010_0_x_00;
      patterns[1166] = 32'b0101001001000000_1_xx_100_xxx_010_0_1_01;
      patterns[1167] = 32'b0100001001000000_0_xx_100_010_xxx_1_x_xx;
      patterns[1168] = 32'b0000001010001100_1_xx_xxx_xxx_010_0_x_10;
      patterns[1169] = 32'b1000001001000111_1_00_100_111_010_0_x_00;
      patterns[1170] = 32'b1001001001000111_1_01_100_111_010_0_x_00;
      patterns[1171] = 32'b1010001001000111_1_10_100_111_010_0_x_00;
      patterns[1172] = 32'b1011001001000111_1_11_100_111_010_0_x_00;
      patterns[1173] = 32'b0101001001000000_1_xx_100_xxx_010_0_1_01;
      patterns[1174] = 32'b0100001001000000_0_xx_100_010_xxx_1_x_xx;
      patterns[1175] = 32'b0000001010010101_1_xx_xxx_xxx_010_0_x_10;
      patterns[1176] = 32'b1000001001010000_1_00_101_000_010_0_x_00;
      patterns[1177] = 32'b1001001001010000_1_01_101_000_010_0_x_00;
      patterns[1178] = 32'b1010001001010000_1_10_101_000_010_0_x_00;
      patterns[1179] = 32'b1011001001010000_1_11_101_000_010_0_x_00;
      patterns[1180] = 32'b0101001001010000_1_xx_101_xxx_010_0_1_01;
      patterns[1181] = 32'b0100001001010000_0_xx_101_010_xxx_1_x_xx;
      patterns[1182] = 32'b0000001011010001_1_xx_xxx_xxx_010_0_x_10;
      patterns[1183] = 32'b1000001001010001_1_00_101_001_010_0_x_00;
      patterns[1184] = 32'b1001001001010001_1_01_101_001_010_0_x_00;
      patterns[1185] = 32'b1010001001010001_1_10_101_001_010_0_x_00;
      patterns[1186] = 32'b1011001001010001_1_11_101_001_010_0_x_00;
      patterns[1187] = 32'b0101001001010000_1_xx_101_xxx_010_0_1_01;
      patterns[1188] = 32'b0100001001010000_0_xx_101_010_xxx_1_x_xx;
      patterns[1189] = 32'b0000001010101111_1_xx_xxx_xxx_010_0_x_10;
      patterns[1190] = 32'b1000001001010010_1_00_101_010_010_0_x_00;
      patterns[1191] = 32'b1001001001010010_1_01_101_010_010_0_x_00;
      patterns[1192] = 32'b1010001001010010_1_10_101_010_010_0_x_00;
      patterns[1193] = 32'b1011001001010010_1_11_101_010_010_0_x_00;
      patterns[1194] = 32'b0101001001010000_1_xx_101_xxx_010_0_1_01;
      patterns[1195] = 32'b0100001001010000_0_xx_101_010_xxx_1_x_xx;
      patterns[1196] = 32'b0000001011001001_1_xx_xxx_xxx_010_0_x_10;
      patterns[1197] = 32'b1000001001010011_1_00_101_011_010_0_x_00;
      patterns[1198] = 32'b1001001001010011_1_01_101_011_010_0_x_00;
      patterns[1199] = 32'b1010001001010011_1_10_101_011_010_0_x_00;
      patterns[1200] = 32'b1011001001010011_1_11_101_011_010_0_x_00;
      patterns[1201] = 32'b0101001001010000_1_xx_101_xxx_010_0_1_01;
      patterns[1202] = 32'b0100001001010000_0_xx_101_010_xxx_1_x_xx;
      patterns[1203] = 32'b0000001001100111_1_xx_xxx_xxx_010_0_x_10;
      patterns[1204] = 32'b1000001001010100_1_00_101_100_010_0_x_00;
      patterns[1205] = 32'b1001001001010100_1_01_101_100_010_0_x_00;
      patterns[1206] = 32'b1010001001010100_1_10_101_100_010_0_x_00;
      patterns[1207] = 32'b1011001001010100_1_11_101_100_010_0_x_00;
      patterns[1208] = 32'b0101001001010000_1_xx_101_xxx_010_0_1_01;
      patterns[1209] = 32'b0100001001010000_0_xx_101_010_xxx_1_x_xx;
      patterns[1210] = 32'b0000001001111011_1_xx_xxx_xxx_010_0_x_10;
      patterns[1211] = 32'b1000001001010101_1_00_101_101_010_0_x_00;
      patterns[1212] = 32'b1001001001010101_1_01_101_101_010_0_x_00;
      patterns[1213] = 32'b1010001001010101_1_10_101_101_010_0_x_00;
      patterns[1214] = 32'b1011001001010101_1_11_101_101_010_0_x_00;
      patterns[1215] = 32'b0101001001010000_1_xx_101_xxx_010_0_1_01;
      patterns[1216] = 32'b0100001001010000_0_xx_101_010_xxx_1_x_xx;
      patterns[1217] = 32'b0000001001000010_1_xx_xxx_xxx_010_0_x_10;
      patterns[1218] = 32'b1000001001010110_1_00_101_110_010_0_x_00;
      patterns[1219] = 32'b1001001001010110_1_01_101_110_010_0_x_00;
      patterns[1220] = 32'b1010001001010110_1_10_101_110_010_0_x_00;
      patterns[1221] = 32'b1011001001010110_1_11_101_110_010_0_x_00;
      patterns[1222] = 32'b0101001001010000_1_xx_101_xxx_010_0_1_01;
      patterns[1223] = 32'b0100001001010000_0_xx_101_010_xxx_1_x_xx;
      patterns[1224] = 32'b0000001010011110_1_xx_xxx_xxx_010_0_x_10;
      patterns[1225] = 32'b1000001001010111_1_00_101_111_010_0_x_00;
      patterns[1226] = 32'b1001001001010111_1_01_101_111_010_0_x_00;
      patterns[1227] = 32'b1010001001010111_1_10_101_111_010_0_x_00;
      patterns[1228] = 32'b1011001001010111_1_11_101_111_010_0_x_00;
      patterns[1229] = 32'b0101001001010000_1_xx_101_xxx_010_0_1_01;
      patterns[1230] = 32'b0100001001010000_0_xx_101_010_xxx_1_x_xx;
      patterns[1231] = 32'b0000001000000001_1_xx_xxx_xxx_010_0_x_10;
      patterns[1232] = 32'b1000001001100000_1_00_110_000_010_0_x_00;
      patterns[1233] = 32'b1001001001100000_1_01_110_000_010_0_x_00;
      patterns[1234] = 32'b1010001001100000_1_10_110_000_010_0_x_00;
      patterns[1235] = 32'b1011001001100000_1_11_110_000_010_0_x_00;
      patterns[1236] = 32'b0101001001100000_1_xx_110_xxx_010_0_1_01;
      patterns[1237] = 32'b0100001001100000_0_xx_110_010_xxx_1_x_xx;
      patterns[1238] = 32'b0000001000001110_1_xx_xxx_xxx_010_0_x_10;
      patterns[1239] = 32'b1000001001100001_1_00_110_001_010_0_x_00;
      patterns[1240] = 32'b1001001001100001_1_01_110_001_010_0_x_00;
      patterns[1241] = 32'b1010001001100001_1_10_110_001_010_0_x_00;
      patterns[1242] = 32'b1011001001100001_1_11_110_001_010_0_x_00;
      patterns[1243] = 32'b0101001001100000_1_xx_110_xxx_010_0_1_01;
      patterns[1244] = 32'b0100001001100000_0_xx_110_010_xxx_1_x_xx;
      patterns[1245] = 32'b0000001000011111_1_xx_xxx_xxx_010_0_x_10;
      patterns[1246] = 32'b1000001001100010_1_00_110_010_010_0_x_00;
      patterns[1247] = 32'b1001001001100010_1_01_110_010_010_0_x_00;
      patterns[1248] = 32'b1010001001100010_1_10_110_010_010_0_x_00;
      patterns[1249] = 32'b1011001001100010_1_11_110_010_010_0_x_00;
      patterns[1250] = 32'b0101001001100000_1_xx_110_xxx_010_0_1_01;
      patterns[1251] = 32'b0100001001100000_0_xx_110_010_xxx_1_x_xx;
      patterns[1252] = 32'b0000001001110000_1_xx_xxx_xxx_010_0_x_10;
      patterns[1253] = 32'b1000001001100011_1_00_110_011_010_0_x_00;
      patterns[1254] = 32'b1001001001100011_1_01_110_011_010_0_x_00;
      patterns[1255] = 32'b1010001001100011_1_10_110_011_010_0_x_00;
      patterns[1256] = 32'b1011001001100011_1_11_110_011_010_0_x_00;
      patterns[1257] = 32'b0101001001100000_1_xx_110_xxx_010_0_1_01;
      patterns[1258] = 32'b0100001001100000_0_xx_110_010_xxx_1_x_xx;
      patterns[1259] = 32'b0000001011110010_1_xx_xxx_xxx_010_0_x_10;
      patterns[1260] = 32'b1000001001100100_1_00_110_100_010_0_x_00;
      patterns[1261] = 32'b1001001001100100_1_01_110_100_010_0_x_00;
      patterns[1262] = 32'b1010001001100100_1_10_110_100_010_0_x_00;
      patterns[1263] = 32'b1011001001100100_1_11_110_100_010_0_x_00;
      patterns[1264] = 32'b0101001001100000_1_xx_110_xxx_010_0_1_01;
      patterns[1265] = 32'b0100001001100000_0_xx_110_010_xxx_1_x_xx;
      patterns[1266] = 32'b0000001001100001_1_xx_xxx_xxx_010_0_x_10;
      patterns[1267] = 32'b1000001001100101_1_00_110_101_010_0_x_00;
      patterns[1268] = 32'b1001001001100101_1_01_110_101_010_0_x_00;
      patterns[1269] = 32'b1010001001100101_1_10_110_101_010_0_x_00;
      patterns[1270] = 32'b1011001001100101_1_11_110_101_010_0_x_00;
      patterns[1271] = 32'b0101001001100000_1_xx_110_xxx_010_0_1_01;
      patterns[1272] = 32'b0100001001100000_0_xx_110_010_xxx_1_x_xx;
      patterns[1273] = 32'b0000001011100000_1_xx_xxx_xxx_010_0_x_10;
      patterns[1274] = 32'b1000001001100110_1_00_110_110_010_0_x_00;
      patterns[1275] = 32'b1001001001100110_1_01_110_110_010_0_x_00;
      patterns[1276] = 32'b1010001001100110_1_10_110_110_010_0_x_00;
      patterns[1277] = 32'b1011001001100110_1_11_110_110_010_0_x_00;
      patterns[1278] = 32'b0101001001100000_1_xx_110_xxx_010_0_1_01;
      patterns[1279] = 32'b0100001001100000_0_xx_110_010_xxx_1_x_xx;
      patterns[1280] = 32'b0000001000100000_1_xx_xxx_xxx_010_0_x_10;
      patterns[1281] = 32'b1000001001100111_1_00_110_111_010_0_x_00;
      patterns[1282] = 32'b1001001001100111_1_01_110_111_010_0_x_00;
      patterns[1283] = 32'b1010001001100111_1_10_110_111_010_0_x_00;
      patterns[1284] = 32'b1011001001100111_1_11_110_111_010_0_x_00;
      patterns[1285] = 32'b0101001001100000_1_xx_110_xxx_010_0_1_01;
      patterns[1286] = 32'b0100001001100000_0_xx_110_010_xxx_1_x_xx;
      patterns[1287] = 32'b0000001000011100_1_xx_xxx_xxx_010_0_x_10;
      patterns[1288] = 32'b1000001001110000_1_00_111_000_010_0_x_00;
      patterns[1289] = 32'b1001001001110000_1_01_111_000_010_0_x_00;
      patterns[1290] = 32'b1010001001110000_1_10_111_000_010_0_x_00;
      patterns[1291] = 32'b1011001001110000_1_11_111_000_010_0_x_00;
      patterns[1292] = 32'b0101001001110000_1_xx_111_xxx_010_0_1_01;
      patterns[1293] = 32'b0100001001110000_0_xx_111_010_xxx_1_x_xx;
      patterns[1294] = 32'b0000001010110011_1_xx_xxx_xxx_010_0_x_10;
      patterns[1295] = 32'b1000001001110001_1_00_111_001_010_0_x_00;
      patterns[1296] = 32'b1001001001110001_1_01_111_001_010_0_x_00;
      patterns[1297] = 32'b1010001001110001_1_10_111_001_010_0_x_00;
      patterns[1298] = 32'b1011001001110001_1_11_111_001_010_0_x_00;
      patterns[1299] = 32'b0101001001110000_1_xx_111_xxx_010_0_1_01;
      patterns[1300] = 32'b0100001001110000_0_xx_111_010_xxx_1_x_xx;
      patterns[1301] = 32'b0000001010000100_1_xx_xxx_xxx_010_0_x_10;
      patterns[1302] = 32'b1000001001110010_1_00_111_010_010_0_x_00;
      patterns[1303] = 32'b1001001001110010_1_01_111_010_010_0_x_00;
      patterns[1304] = 32'b1010001001110010_1_10_111_010_010_0_x_00;
      patterns[1305] = 32'b1011001001110010_1_11_111_010_010_0_x_00;
      patterns[1306] = 32'b0101001001110000_1_xx_111_xxx_010_0_1_01;
      patterns[1307] = 32'b0100001001110000_0_xx_111_010_xxx_1_x_xx;
      patterns[1308] = 32'b0000001001000010_1_xx_xxx_xxx_010_0_x_10;
      patterns[1309] = 32'b1000001001110011_1_00_111_011_010_0_x_00;
      patterns[1310] = 32'b1001001001110011_1_01_111_011_010_0_x_00;
      patterns[1311] = 32'b1010001001110011_1_10_111_011_010_0_x_00;
      patterns[1312] = 32'b1011001001110011_1_11_111_011_010_0_x_00;
      patterns[1313] = 32'b0101001001110000_1_xx_111_xxx_010_0_1_01;
      patterns[1314] = 32'b0100001001110000_0_xx_111_010_xxx_1_x_xx;
      patterns[1315] = 32'b0000001011110101_1_xx_xxx_xxx_010_0_x_10;
      patterns[1316] = 32'b1000001001110100_1_00_111_100_010_0_x_00;
      patterns[1317] = 32'b1001001001110100_1_01_111_100_010_0_x_00;
      patterns[1318] = 32'b1010001001110100_1_10_111_100_010_0_x_00;
      patterns[1319] = 32'b1011001001110100_1_11_111_100_010_0_x_00;
      patterns[1320] = 32'b0101001001110000_1_xx_111_xxx_010_0_1_01;
      patterns[1321] = 32'b0100001001110000_0_xx_111_010_xxx_1_x_xx;
      patterns[1322] = 32'b0000001001000001_1_xx_xxx_xxx_010_0_x_10;
      patterns[1323] = 32'b1000001001110101_1_00_111_101_010_0_x_00;
      patterns[1324] = 32'b1001001001110101_1_01_111_101_010_0_x_00;
      patterns[1325] = 32'b1010001001110101_1_10_111_101_010_0_x_00;
      patterns[1326] = 32'b1011001001110101_1_11_111_101_010_0_x_00;
      patterns[1327] = 32'b0101001001110000_1_xx_111_xxx_010_0_1_01;
      patterns[1328] = 32'b0100001001110000_0_xx_111_010_xxx_1_x_xx;
      patterns[1329] = 32'b0000001010000110_1_xx_xxx_xxx_010_0_x_10;
      patterns[1330] = 32'b1000001001110110_1_00_111_110_010_0_x_00;
      patterns[1331] = 32'b1001001001110110_1_01_111_110_010_0_x_00;
      patterns[1332] = 32'b1010001001110110_1_10_111_110_010_0_x_00;
      patterns[1333] = 32'b1011001001110110_1_11_111_110_010_0_x_00;
      patterns[1334] = 32'b0101001001110000_1_xx_111_xxx_010_0_1_01;
      patterns[1335] = 32'b0100001001110000_0_xx_111_010_xxx_1_x_xx;
      patterns[1336] = 32'b0000001010110010_1_xx_xxx_xxx_010_0_x_10;
      patterns[1337] = 32'b1000001001110111_1_00_111_111_010_0_x_00;
      patterns[1338] = 32'b1001001001110111_1_01_111_111_010_0_x_00;
      patterns[1339] = 32'b1010001001110111_1_10_111_111_010_0_x_00;
      patterns[1340] = 32'b1011001001110111_1_11_111_111_010_0_x_00;
      patterns[1341] = 32'b0101001001110000_1_xx_111_xxx_010_0_1_01;
      patterns[1342] = 32'b0100001001110000_0_xx_111_010_xxx_1_x_xx;
      patterns[1343] = 32'b0000001010000000_1_xx_xxx_xxx_010_0_x_10;
      patterns[1344] = 32'b1000001100000000_1_00_000_000_011_0_x_00;
      patterns[1345] = 32'b1001001100000000_1_01_000_000_011_0_x_00;
      patterns[1346] = 32'b1010001100000000_1_10_000_000_011_0_x_00;
      patterns[1347] = 32'b1011001100000000_1_11_000_000_011_0_x_00;
      patterns[1348] = 32'b0101001100000000_1_xx_000_xxx_011_0_1_01;
      patterns[1349] = 32'b0100001100000000_0_xx_000_011_xxx_1_x_xx;
      patterns[1350] = 32'b0000001100010011_1_xx_xxx_xxx_011_0_x_10;
      patterns[1351] = 32'b1000001100000001_1_00_000_001_011_0_x_00;
      patterns[1352] = 32'b1001001100000001_1_01_000_001_011_0_x_00;
      patterns[1353] = 32'b1010001100000001_1_10_000_001_011_0_x_00;
      patterns[1354] = 32'b1011001100000001_1_11_000_001_011_0_x_00;
      patterns[1355] = 32'b0101001100000000_1_xx_000_xxx_011_0_1_01;
      patterns[1356] = 32'b0100001100000000_0_xx_000_011_xxx_1_x_xx;
      patterns[1357] = 32'b0000001101011100_1_xx_xxx_xxx_011_0_x_10;
      patterns[1358] = 32'b1000001100000010_1_00_000_010_011_0_x_00;
      patterns[1359] = 32'b1001001100000010_1_01_000_010_011_0_x_00;
      patterns[1360] = 32'b1010001100000010_1_10_000_010_011_0_x_00;
      patterns[1361] = 32'b1011001100000010_1_11_000_010_011_0_x_00;
      patterns[1362] = 32'b0101001100000000_1_xx_000_xxx_011_0_1_01;
      patterns[1363] = 32'b0100001100000000_0_xx_000_011_xxx_1_x_xx;
      patterns[1364] = 32'b0000001110101000_1_xx_xxx_xxx_011_0_x_10;
      patterns[1365] = 32'b1000001100000011_1_00_000_011_011_0_x_00;
      patterns[1366] = 32'b1001001100000011_1_01_000_011_011_0_x_00;
      patterns[1367] = 32'b1010001100000011_1_10_000_011_011_0_x_00;
      patterns[1368] = 32'b1011001100000011_1_11_000_011_011_0_x_00;
      patterns[1369] = 32'b0101001100000000_1_xx_000_xxx_011_0_1_01;
      patterns[1370] = 32'b0100001100000000_0_xx_000_011_xxx_1_x_xx;
      patterns[1371] = 32'b0000001100001010_1_xx_xxx_xxx_011_0_x_10;
      patterns[1372] = 32'b1000001100000100_1_00_000_100_011_0_x_00;
      patterns[1373] = 32'b1001001100000100_1_01_000_100_011_0_x_00;
      patterns[1374] = 32'b1010001100000100_1_10_000_100_011_0_x_00;
      patterns[1375] = 32'b1011001100000100_1_11_000_100_011_0_x_00;
      patterns[1376] = 32'b0101001100000000_1_xx_000_xxx_011_0_1_01;
      patterns[1377] = 32'b0100001100000000_0_xx_000_011_xxx_1_x_xx;
      patterns[1378] = 32'b0000001110111100_1_xx_xxx_xxx_011_0_x_10;
      patterns[1379] = 32'b1000001100000101_1_00_000_101_011_0_x_00;
      patterns[1380] = 32'b1001001100000101_1_01_000_101_011_0_x_00;
      patterns[1381] = 32'b1010001100000101_1_10_000_101_011_0_x_00;
      patterns[1382] = 32'b1011001100000101_1_11_000_101_011_0_x_00;
      patterns[1383] = 32'b0101001100000000_1_xx_000_xxx_011_0_1_01;
      patterns[1384] = 32'b0100001100000000_0_xx_000_011_xxx_1_x_xx;
      patterns[1385] = 32'b0000001101000111_1_xx_xxx_xxx_011_0_x_10;
      patterns[1386] = 32'b1000001100000110_1_00_000_110_011_0_x_00;
      patterns[1387] = 32'b1001001100000110_1_01_000_110_011_0_x_00;
      patterns[1388] = 32'b1010001100000110_1_10_000_110_011_0_x_00;
      patterns[1389] = 32'b1011001100000110_1_11_000_110_011_0_x_00;
      patterns[1390] = 32'b0101001100000000_1_xx_000_xxx_011_0_1_01;
      patterns[1391] = 32'b0100001100000000_0_xx_000_011_xxx_1_x_xx;
      patterns[1392] = 32'b0000001100000101_1_xx_xxx_xxx_011_0_x_10;
      patterns[1393] = 32'b1000001100000111_1_00_000_111_011_0_x_00;
      patterns[1394] = 32'b1001001100000111_1_01_000_111_011_0_x_00;
      patterns[1395] = 32'b1010001100000111_1_10_000_111_011_0_x_00;
      patterns[1396] = 32'b1011001100000111_1_11_000_111_011_0_x_00;
      patterns[1397] = 32'b0101001100000000_1_xx_000_xxx_011_0_1_01;
      patterns[1398] = 32'b0100001100000000_0_xx_000_011_xxx_1_x_xx;
      patterns[1399] = 32'b0000001111011011_1_xx_xxx_xxx_011_0_x_10;
      patterns[1400] = 32'b1000001100010000_1_00_001_000_011_0_x_00;
      patterns[1401] = 32'b1001001100010000_1_01_001_000_011_0_x_00;
      patterns[1402] = 32'b1010001100010000_1_10_001_000_011_0_x_00;
      patterns[1403] = 32'b1011001100010000_1_11_001_000_011_0_x_00;
      patterns[1404] = 32'b0101001100010000_1_xx_001_xxx_011_0_1_01;
      patterns[1405] = 32'b0100001100010000_0_xx_001_011_xxx_1_x_xx;
      patterns[1406] = 32'b0000001111000000_1_xx_xxx_xxx_011_0_x_10;
      patterns[1407] = 32'b1000001100010001_1_00_001_001_011_0_x_00;
      patterns[1408] = 32'b1001001100010001_1_01_001_001_011_0_x_00;
      patterns[1409] = 32'b1010001100010001_1_10_001_001_011_0_x_00;
      patterns[1410] = 32'b1011001100010001_1_11_001_001_011_0_x_00;
      patterns[1411] = 32'b0101001100010000_1_xx_001_xxx_011_0_1_01;
      patterns[1412] = 32'b0100001100010000_0_xx_001_011_xxx_1_x_xx;
      patterns[1413] = 32'b0000001111011001_1_xx_xxx_xxx_011_0_x_10;
      patterns[1414] = 32'b1000001100010010_1_00_001_010_011_0_x_00;
      patterns[1415] = 32'b1001001100010010_1_01_001_010_011_0_x_00;
      patterns[1416] = 32'b1010001100010010_1_10_001_010_011_0_x_00;
      patterns[1417] = 32'b1011001100010010_1_11_001_010_011_0_x_00;
      patterns[1418] = 32'b0101001100010000_1_xx_001_xxx_011_0_1_01;
      patterns[1419] = 32'b0100001100010000_0_xx_001_011_xxx_1_x_xx;
      patterns[1420] = 32'b0000001111101001_1_xx_xxx_xxx_011_0_x_10;
      patterns[1421] = 32'b1000001100010011_1_00_001_011_011_0_x_00;
      patterns[1422] = 32'b1001001100010011_1_01_001_011_011_0_x_00;
      patterns[1423] = 32'b1010001100010011_1_10_001_011_011_0_x_00;
      patterns[1424] = 32'b1011001100010011_1_11_001_011_011_0_x_00;
      patterns[1425] = 32'b0101001100010000_1_xx_001_xxx_011_0_1_01;
      patterns[1426] = 32'b0100001100010000_0_xx_001_011_xxx_1_x_xx;
      patterns[1427] = 32'b0000001111110010_1_xx_xxx_xxx_011_0_x_10;
      patterns[1428] = 32'b1000001100010100_1_00_001_100_011_0_x_00;
      patterns[1429] = 32'b1001001100010100_1_01_001_100_011_0_x_00;
      patterns[1430] = 32'b1010001100010100_1_10_001_100_011_0_x_00;
      patterns[1431] = 32'b1011001100010100_1_11_001_100_011_0_x_00;
      patterns[1432] = 32'b0101001100010000_1_xx_001_xxx_011_0_1_01;
      patterns[1433] = 32'b0100001100010000_0_xx_001_011_xxx_1_x_xx;
      patterns[1434] = 32'b0000001100101101_1_xx_xxx_xxx_011_0_x_10;
      patterns[1435] = 32'b1000001100010101_1_00_001_101_011_0_x_00;
      patterns[1436] = 32'b1001001100010101_1_01_001_101_011_0_x_00;
      patterns[1437] = 32'b1010001100010101_1_10_001_101_011_0_x_00;
      patterns[1438] = 32'b1011001100010101_1_11_001_101_011_0_x_00;
      patterns[1439] = 32'b0101001100010000_1_xx_001_xxx_011_0_1_01;
      patterns[1440] = 32'b0100001100010000_0_xx_001_011_xxx_1_x_xx;
      patterns[1441] = 32'b0000001101010100_1_xx_xxx_xxx_011_0_x_10;
      patterns[1442] = 32'b1000001100010110_1_00_001_110_011_0_x_00;
      patterns[1443] = 32'b1001001100010110_1_01_001_110_011_0_x_00;
      patterns[1444] = 32'b1010001100010110_1_10_001_110_011_0_x_00;
      patterns[1445] = 32'b1011001100010110_1_11_001_110_011_0_x_00;
      patterns[1446] = 32'b0101001100010000_1_xx_001_xxx_011_0_1_01;
      patterns[1447] = 32'b0100001100010000_0_xx_001_011_xxx_1_x_xx;
      patterns[1448] = 32'b0000001110011001_1_xx_xxx_xxx_011_0_x_10;
      patterns[1449] = 32'b1000001100010111_1_00_001_111_011_0_x_00;
      patterns[1450] = 32'b1001001100010111_1_01_001_111_011_0_x_00;
      patterns[1451] = 32'b1010001100010111_1_10_001_111_011_0_x_00;
      patterns[1452] = 32'b1011001100010111_1_11_001_111_011_0_x_00;
      patterns[1453] = 32'b0101001100010000_1_xx_001_xxx_011_0_1_01;
      patterns[1454] = 32'b0100001100010000_0_xx_001_011_xxx_1_x_xx;
      patterns[1455] = 32'b0000001111101000_1_xx_xxx_xxx_011_0_x_10;
      patterns[1456] = 32'b1000001100100000_1_00_010_000_011_0_x_00;
      patterns[1457] = 32'b1001001100100000_1_01_010_000_011_0_x_00;
      patterns[1458] = 32'b1010001100100000_1_10_010_000_011_0_x_00;
      patterns[1459] = 32'b1011001100100000_1_11_010_000_011_0_x_00;
      patterns[1460] = 32'b0101001100100000_1_xx_010_xxx_011_0_1_01;
      patterns[1461] = 32'b0100001100100000_0_xx_010_011_xxx_1_x_xx;
      patterns[1462] = 32'b0000001101001110_1_xx_xxx_xxx_011_0_x_10;
      patterns[1463] = 32'b1000001100100001_1_00_010_001_011_0_x_00;
      patterns[1464] = 32'b1001001100100001_1_01_010_001_011_0_x_00;
      patterns[1465] = 32'b1010001100100001_1_10_010_001_011_0_x_00;
      patterns[1466] = 32'b1011001100100001_1_11_010_001_011_0_x_00;
      patterns[1467] = 32'b0101001100100000_1_xx_010_xxx_011_0_1_01;
      patterns[1468] = 32'b0100001100100000_0_xx_010_011_xxx_1_x_xx;
      patterns[1469] = 32'b0000001101001110_1_xx_xxx_xxx_011_0_x_10;
      patterns[1470] = 32'b1000001100100010_1_00_010_010_011_0_x_00;
      patterns[1471] = 32'b1001001100100010_1_01_010_010_011_0_x_00;
      patterns[1472] = 32'b1010001100100010_1_10_010_010_011_0_x_00;
      patterns[1473] = 32'b1011001100100010_1_11_010_010_011_0_x_00;
      patterns[1474] = 32'b0101001100100000_1_xx_010_xxx_011_0_1_01;
      patterns[1475] = 32'b0100001100100000_0_xx_010_011_xxx_1_x_xx;
      patterns[1476] = 32'b0000001101010001_1_xx_xxx_xxx_011_0_x_10;
      patterns[1477] = 32'b1000001100100011_1_00_010_011_011_0_x_00;
      patterns[1478] = 32'b1001001100100011_1_01_010_011_011_0_x_00;
      patterns[1479] = 32'b1010001100100011_1_10_010_011_011_0_x_00;
      patterns[1480] = 32'b1011001100100011_1_11_010_011_011_0_x_00;
      patterns[1481] = 32'b0101001100100000_1_xx_010_xxx_011_0_1_01;
      patterns[1482] = 32'b0100001100100000_0_xx_010_011_xxx_1_x_xx;
      patterns[1483] = 32'b0000001111001110_1_xx_xxx_xxx_011_0_x_10;
      patterns[1484] = 32'b1000001100100100_1_00_010_100_011_0_x_00;
      patterns[1485] = 32'b1001001100100100_1_01_010_100_011_0_x_00;
      patterns[1486] = 32'b1010001100100100_1_10_010_100_011_0_x_00;
      patterns[1487] = 32'b1011001100100100_1_11_010_100_011_0_x_00;
      patterns[1488] = 32'b0101001100100000_1_xx_010_xxx_011_0_1_01;
      patterns[1489] = 32'b0100001100100000_0_xx_010_011_xxx_1_x_xx;
      patterns[1490] = 32'b0000001110001110_1_xx_xxx_xxx_011_0_x_10;
      patterns[1491] = 32'b1000001100100101_1_00_010_101_011_0_x_00;
      patterns[1492] = 32'b1001001100100101_1_01_010_101_011_0_x_00;
      patterns[1493] = 32'b1010001100100101_1_10_010_101_011_0_x_00;
      patterns[1494] = 32'b1011001100100101_1_11_010_101_011_0_x_00;
      patterns[1495] = 32'b0101001100100000_1_xx_010_xxx_011_0_1_01;
      patterns[1496] = 32'b0100001100100000_0_xx_010_011_xxx_1_x_xx;
      patterns[1497] = 32'b0000001110110000_1_xx_xxx_xxx_011_0_x_10;
      patterns[1498] = 32'b1000001100100110_1_00_010_110_011_0_x_00;
      patterns[1499] = 32'b1001001100100110_1_01_010_110_011_0_x_00;
      patterns[1500] = 32'b1010001100100110_1_10_010_110_011_0_x_00;
      patterns[1501] = 32'b1011001100100110_1_11_010_110_011_0_x_00;
      patterns[1502] = 32'b0101001100100000_1_xx_010_xxx_011_0_1_01;
      patterns[1503] = 32'b0100001100100000_0_xx_010_011_xxx_1_x_xx;
      patterns[1504] = 32'b0000001100000001_1_xx_xxx_xxx_011_0_x_10;
      patterns[1505] = 32'b1000001100100111_1_00_010_111_011_0_x_00;
      patterns[1506] = 32'b1001001100100111_1_01_010_111_011_0_x_00;
      patterns[1507] = 32'b1010001100100111_1_10_010_111_011_0_x_00;
      patterns[1508] = 32'b1011001100100111_1_11_010_111_011_0_x_00;
      patterns[1509] = 32'b0101001100100000_1_xx_010_xxx_011_0_1_01;
      patterns[1510] = 32'b0100001100100000_0_xx_010_011_xxx_1_x_xx;
      patterns[1511] = 32'b0000001110101111_1_xx_xxx_xxx_011_0_x_10;
      patterns[1512] = 32'b1000001100110000_1_00_011_000_011_0_x_00;
      patterns[1513] = 32'b1001001100110000_1_01_011_000_011_0_x_00;
      patterns[1514] = 32'b1010001100110000_1_10_011_000_011_0_x_00;
      patterns[1515] = 32'b1011001100110000_1_11_011_000_011_0_x_00;
      patterns[1516] = 32'b0101001100110000_1_xx_011_xxx_011_0_1_01;
      patterns[1517] = 32'b0100001100110000_0_xx_011_011_xxx_1_x_xx;
      patterns[1518] = 32'b0000001100100111_1_xx_xxx_xxx_011_0_x_10;
      patterns[1519] = 32'b1000001100110001_1_00_011_001_011_0_x_00;
      patterns[1520] = 32'b1001001100110001_1_01_011_001_011_0_x_00;
      patterns[1521] = 32'b1010001100110001_1_10_011_001_011_0_x_00;
      patterns[1522] = 32'b1011001100110001_1_11_011_001_011_0_x_00;
      patterns[1523] = 32'b0101001100110000_1_xx_011_xxx_011_0_1_01;
      patterns[1524] = 32'b0100001100110000_0_xx_011_011_xxx_1_x_xx;
      patterns[1525] = 32'b0000001100101000_1_xx_xxx_xxx_011_0_x_10;
      patterns[1526] = 32'b1000001100110010_1_00_011_010_011_0_x_00;
      patterns[1527] = 32'b1001001100110010_1_01_011_010_011_0_x_00;
      patterns[1528] = 32'b1010001100110010_1_10_011_010_011_0_x_00;
      patterns[1529] = 32'b1011001100110010_1_11_011_010_011_0_x_00;
      patterns[1530] = 32'b0101001100110000_1_xx_011_xxx_011_0_1_01;
      patterns[1531] = 32'b0100001100110000_0_xx_011_011_xxx_1_x_xx;
      patterns[1532] = 32'b0000001110110001_1_xx_xxx_xxx_011_0_x_10;
      patterns[1533] = 32'b1000001100110011_1_00_011_011_011_0_x_00;
      patterns[1534] = 32'b1001001100110011_1_01_011_011_011_0_x_00;
      patterns[1535] = 32'b1010001100110011_1_10_011_011_011_0_x_00;
      patterns[1536] = 32'b1011001100110011_1_11_011_011_011_0_x_00;
      patterns[1537] = 32'b0101001100110000_1_xx_011_xxx_011_0_1_01;
      patterns[1538] = 32'b0100001100110000_0_xx_011_011_xxx_1_x_xx;
      patterns[1539] = 32'b0000001111100001_1_xx_xxx_xxx_011_0_x_10;
      patterns[1540] = 32'b1000001100110100_1_00_011_100_011_0_x_00;
      patterns[1541] = 32'b1001001100110100_1_01_011_100_011_0_x_00;
      patterns[1542] = 32'b1010001100110100_1_10_011_100_011_0_x_00;
      patterns[1543] = 32'b1011001100110100_1_11_011_100_011_0_x_00;
      patterns[1544] = 32'b0101001100110000_1_xx_011_xxx_011_0_1_01;
      patterns[1545] = 32'b0100001100110000_0_xx_011_011_xxx_1_x_xx;
      patterns[1546] = 32'b0000001111101110_1_xx_xxx_xxx_011_0_x_10;
      patterns[1547] = 32'b1000001100110101_1_00_011_101_011_0_x_00;
      patterns[1548] = 32'b1001001100110101_1_01_011_101_011_0_x_00;
      patterns[1549] = 32'b1010001100110101_1_10_011_101_011_0_x_00;
      patterns[1550] = 32'b1011001100110101_1_11_011_101_011_0_x_00;
      patterns[1551] = 32'b0101001100110000_1_xx_011_xxx_011_0_1_01;
      patterns[1552] = 32'b0100001100110000_0_xx_011_011_xxx_1_x_xx;
      patterns[1553] = 32'b0000001110100000_1_xx_xxx_xxx_011_0_x_10;
      patterns[1554] = 32'b1000001100110110_1_00_011_110_011_0_x_00;
      patterns[1555] = 32'b1001001100110110_1_01_011_110_011_0_x_00;
      patterns[1556] = 32'b1010001100110110_1_10_011_110_011_0_x_00;
      patterns[1557] = 32'b1011001100110110_1_11_011_110_011_0_x_00;
      patterns[1558] = 32'b0101001100110000_1_xx_011_xxx_011_0_1_01;
      patterns[1559] = 32'b0100001100110000_0_xx_011_011_xxx_1_x_xx;
      patterns[1560] = 32'b0000001100100011_1_xx_xxx_xxx_011_0_x_10;
      patterns[1561] = 32'b1000001100110111_1_00_011_111_011_0_x_00;
      patterns[1562] = 32'b1001001100110111_1_01_011_111_011_0_x_00;
      patterns[1563] = 32'b1010001100110111_1_10_011_111_011_0_x_00;
      patterns[1564] = 32'b1011001100110111_1_11_011_111_011_0_x_00;
      patterns[1565] = 32'b0101001100110000_1_xx_011_xxx_011_0_1_01;
      patterns[1566] = 32'b0100001100110000_0_xx_011_011_xxx_1_x_xx;
      patterns[1567] = 32'b0000001111111011_1_xx_xxx_xxx_011_0_x_10;
      patterns[1568] = 32'b1000001101000000_1_00_100_000_011_0_x_00;
      patterns[1569] = 32'b1001001101000000_1_01_100_000_011_0_x_00;
      patterns[1570] = 32'b1010001101000000_1_10_100_000_011_0_x_00;
      patterns[1571] = 32'b1011001101000000_1_11_100_000_011_0_x_00;
      patterns[1572] = 32'b0101001101000000_1_xx_100_xxx_011_0_1_01;
      patterns[1573] = 32'b0100001101000000_0_xx_100_011_xxx_1_x_xx;
      patterns[1574] = 32'b0000001100110111_1_xx_xxx_xxx_011_0_x_10;
      patterns[1575] = 32'b1000001101000001_1_00_100_001_011_0_x_00;
      patterns[1576] = 32'b1001001101000001_1_01_100_001_011_0_x_00;
      patterns[1577] = 32'b1010001101000001_1_10_100_001_011_0_x_00;
      patterns[1578] = 32'b1011001101000001_1_11_100_001_011_0_x_00;
      patterns[1579] = 32'b0101001101000000_1_xx_100_xxx_011_0_1_01;
      patterns[1580] = 32'b0100001101000000_0_xx_100_011_xxx_1_x_xx;
      patterns[1581] = 32'b0000001100110011_1_xx_xxx_xxx_011_0_x_10;
      patterns[1582] = 32'b1000001101000010_1_00_100_010_011_0_x_00;
      patterns[1583] = 32'b1001001101000010_1_01_100_010_011_0_x_00;
      patterns[1584] = 32'b1010001101000010_1_10_100_010_011_0_x_00;
      patterns[1585] = 32'b1011001101000010_1_11_100_010_011_0_x_00;
      patterns[1586] = 32'b0101001101000000_1_xx_100_xxx_011_0_1_01;
      patterns[1587] = 32'b0100001101000000_0_xx_100_011_xxx_1_x_xx;
      patterns[1588] = 32'b0000001101000110_1_xx_xxx_xxx_011_0_x_10;
      patterns[1589] = 32'b1000001101000011_1_00_100_011_011_0_x_00;
      patterns[1590] = 32'b1001001101000011_1_01_100_011_011_0_x_00;
      patterns[1591] = 32'b1010001101000011_1_10_100_011_011_0_x_00;
      patterns[1592] = 32'b1011001101000011_1_11_100_011_011_0_x_00;
      patterns[1593] = 32'b0101001101000000_1_xx_100_xxx_011_0_1_01;
      patterns[1594] = 32'b0100001101000000_0_xx_100_011_xxx_1_x_xx;
      patterns[1595] = 32'b0000001110010001_1_xx_xxx_xxx_011_0_x_10;
      patterns[1596] = 32'b1000001101000100_1_00_100_100_011_0_x_00;
      patterns[1597] = 32'b1001001101000100_1_01_100_100_011_0_x_00;
      patterns[1598] = 32'b1010001101000100_1_10_100_100_011_0_x_00;
      patterns[1599] = 32'b1011001101000100_1_11_100_100_011_0_x_00;
      patterns[1600] = 32'b0101001101000000_1_xx_100_xxx_011_0_1_01;
      patterns[1601] = 32'b0100001101000000_0_xx_100_011_xxx_1_x_xx;
      patterns[1602] = 32'b0000001111011011_1_xx_xxx_xxx_011_0_x_10;
      patterns[1603] = 32'b1000001101000101_1_00_100_101_011_0_x_00;
      patterns[1604] = 32'b1001001101000101_1_01_100_101_011_0_x_00;
      patterns[1605] = 32'b1010001101000101_1_10_100_101_011_0_x_00;
      patterns[1606] = 32'b1011001101000101_1_11_100_101_011_0_x_00;
      patterns[1607] = 32'b0101001101000000_1_xx_100_xxx_011_0_1_01;
      patterns[1608] = 32'b0100001101000000_0_xx_100_011_xxx_1_x_xx;
      patterns[1609] = 32'b0000001101000110_1_xx_xxx_xxx_011_0_x_10;
      patterns[1610] = 32'b1000001101000110_1_00_100_110_011_0_x_00;
      patterns[1611] = 32'b1001001101000110_1_01_100_110_011_0_x_00;
      patterns[1612] = 32'b1010001101000110_1_10_100_110_011_0_x_00;
      patterns[1613] = 32'b1011001101000110_1_11_100_110_011_0_x_00;
      patterns[1614] = 32'b0101001101000000_1_xx_100_xxx_011_0_1_01;
      patterns[1615] = 32'b0100001101000000_0_xx_100_011_xxx_1_x_xx;
      patterns[1616] = 32'b0000001100100010_1_xx_xxx_xxx_011_0_x_10;
      patterns[1617] = 32'b1000001101000111_1_00_100_111_011_0_x_00;
      patterns[1618] = 32'b1001001101000111_1_01_100_111_011_0_x_00;
      patterns[1619] = 32'b1010001101000111_1_10_100_111_011_0_x_00;
      patterns[1620] = 32'b1011001101000111_1_11_100_111_011_0_x_00;
      patterns[1621] = 32'b0101001101000000_1_xx_100_xxx_011_0_1_01;
      patterns[1622] = 32'b0100001101000000_0_xx_100_011_xxx_1_x_xx;
      patterns[1623] = 32'b0000001101011000_1_xx_xxx_xxx_011_0_x_10;
      patterns[1624] = 32'b1000001101010000_1_00_101_000_011_0_x_00;
      patterns[1625] = 32'b1001001101010000_1_01_101_000_011_0_x_00;
      patterns[1626] = 32'b1010001101010000_1_10_101_000_011_0_x_00;
      patterns[1627] = 32'b1011001101010000_1_11_101_000_011_0_x_00;
      patterns[1628] = 32'b0101001101010000_1_xx_101_xxx_011_0_1_01;
      patterns[1629] = 32'b0100001101010000_0_xx_101_011_xxx_1_x_xx;
      patterns[1630] = 32'b0000001101111011_1_xx_xxx_xxx_011_0_x_10;
      patterns[1631] = 32'b1000001101010001_1_00_101_001_011_0_x_00;
      patterns[1632] = 32'b1001001101010001_1_01_101_001_011_0_x_00;
      patterns[1633] = 32'b1010001101010001_1_10_101_001_011_0_x_00;
      patterns[1634] = 32'b1011001101010001_1_11_101_001_011_0_x_00;
      patterns[1635] = 32'b0101001101010000_1_xx_101_xxx_011_0_1_01;
      patterns[1636] = 32'b0100001101010000_0_xx_101_011_xxx_1_x_xx;
      patterns[1637] = 32'b0000001100111100_1_xx_xxx_xxx_011_0_x_10;
      patterns[1638] = 32'b1000001101010010_1_00_101_010_011_0_x_00;
      patterns[1639] = 32'b1001001101010010_1_01_101_010_011_0_x_00;
      patterns[1640] = 32'b1010001101010010_1_10_101_010_011_0_x_00;
      patterns[1641] = 32'b1011001101010010_1_11_101_010_011_0_x_00;
      patterns[1642] = 32'b0101001101010000_1_xx_101_xxx_011_0_1_01;
      patterns[1643] = 32'b0100001101010000_0_xx_101_011_xxx_1_x_xx;
      patterns[1644] = 32'b0000001101100111_1_xx_xxx_xxx_011_0_x_10;
      patterns[1645] = 32'b1000001101010011_1_00_101_011_011_0_x_00;
      patterns[1646] = 32'b1001001101010011_1_01_101_011_011_0_x_00;
      patterns[1647] = 32'b1010001101010011_1_10_101_011_011_0_x_00;
      patterns[1648] = 32'b1011001101010011_1_11_101_011_011_0_x_00;
      patterns[1649] = 32'b0101001101010000_1_xx_101_xxx_011_0_1_01;
      patterns[1650] = 32'b0100001101010000_0_xx_101_011_xxx_1_x_xx;
      patterns[1651] = 32'b0000001101110100_1_xx_xxx_xxx_011_0_x_10;
      patterns[1652] = 32'b1000001101010100_1_00_101_100_011_0_x_00;
      patterns[1653] = 32'b1001001101010100_1_01_101_100_011_0_x_00;
      patterns[1654] = 32'b1010001101010100_1_10_101_100_011_0_x_00;
      patterns[1655] = 32'b1011001101010100_1_11_101_100_011_0_x_00;
      patterns[1656] = 32'b0101001101010000_1_xx_101_xxx_011_0_1_01;
      patterns[1657] = 32'b0100001101010000_0_xx_101_011_xxx_1_x_xx;
      patterns[1658] = 32'b0000001101011110_1_xx_xxx_xxx_011_0_x_10;
      patterns[1659] = 32'b1000001101010101_1_00_101_101_011_0_x_00;
      patterns[1660] = 32'b1001001101010101_1_01_101_101_011_0_x_00;
      patterns[1661] = 32'b1010001101010101_1_10_101_101_011_0_x_00;
      patterns[1662] = 32'b1011001101010101_1_11_101_101_011_0_x_00;
      patterns[1663] = 32'b0101001101010000_1_xx_101_xxx_011_0_1_01;
      patterns[1664] = 32'b0100001101010000_0_xx_101_011_xxx_1_x_xx;
      patterns[1665] = 32'b0000001100100001_1_xx_xxx_xxx_011_0_x_10;
      patterns[1666] = 32'b1000001101010110_1_00_101_110_011_0_x_00;
      patterns[1667] = 32'b1001001101010110_1_01_101_110_011_0_x_00;
      patterns[1668] = 32'b1010001101010110_1_10_101_110_011_0_x_00;
      patterns[1669] = 32'b1011001101010110_1_11_101_110_011_0_x_00;
      patterns[1670] = 32'b0101001101010000_1_xx_101_xxx_011_0_1_01;
      patterns[1671] = 32'b0100001101010000_0_xx_101_011_xxx_1_x_xx;
      patterns[1672] = 32'b0000001111101110_1_xx_xxx_xxx_011_0_x_10;
      patterns[1673] = 32'b1000001101010111_1_00_101_111_011_0_x_00;
      patterns[1674] = 32'b1001001101010111_1_01_101_111_011_0_x_00;
      patterns[1675] = 32'b1010001101010111_1_10_101_111_011_0_x_00;
      patterns[1676] = 32'b1011001101010111_1_11_101_111_011_0_x_00;
      patterns[1677] = 32'b0101001101010000_1_xx_101_xxx_011_0_1_01;
      patterns[1678] = 32'b0100001101010000_0_xx_101_011_xxx_1_x_xx;
      patterns[1679] = 32'b0000001111111001_1_xx_xxx_xxx_011_0_x_10;
      patterns[1680] = 32'b1000001101100000_1_00_110_000_011_0_x_00;
      patterns[1681] = 32'b1001001101100000_1_01_110_000_011_0_x_00;
      patterns[1682] = 32'b1010001101100000_1_10_110_000_011_0_x_00;
      patterns[1683] = 32'b1011001101100000_1_11_110_000_011_0_x_00;
      patterns[1684] = 32'b0101001101100000_1_xx_110_xxx_011_0_1_01;
      patterns[1685] = 32'b0100001101100000_0_xx_110_011_xxx_1_x_xx;
      patterns[1686] = 32'b0000001110101100_1_xx_xxx_xxx_011_0_x_10;
      patterns[1687] = 32'b1000001101100001_1_00_110_001_011_0_x_00;
      patterns[1688] = 32'b1001001101100001_1_01_110_001_011_0_x_00;
      patterns[1689] = 32'b1010001101100001_1_10_110_001_011_0_x_00;
      patterns[1690] = 32'b1011001101100001_1_11_110_001_011_0_x_00;
      patterns[1691] = 32'b0101001101100000_1_xx_110_xxx_011_0_1_01;
      patterns[1692] = 32'b0100001101100000_0_xx_110_011_xxx_1_x_xx;
      patterns[1693] = 32'b0000001101100000_1_xx_xxx_xxx_011_0_x_10;
      patterns[1694] = 32'b1000001101100010_1_00_110_010_011_0_x_00;
      patterns[1695] = 32'b1001001101100010_1_01_110_010_011_0_x_00;
      patterns[1696] = 32'b1010001101100010_1_10_110_010_011_0_x_00;
      patterns[1697] = 32'b1011001101100010_1_11_110_010_011_0_x_00;
      patterns[1698] = 32'b0101001101100000_1_xx_110_xxx_011_0_1_01;
      patterns[1699] = 32'b0100001101100000_0_xx_110_011_xxx_1_x_xx;
      patterns[1700] = 32'b0000001110000100_1_xx_xxx_xxx_011_0_x_10;
      patterns[1701] = 32'b1000001101100011_1_00_110_011_011_0_x_00;
      patterns[1702] = 32'b1001001101100011_1_01_110_011_011_0_x_00;
      patterns[1703] = 32'b1010001101100011_1_10_110_011_011_0_x_00;
      patterns[1704] = 32'b1011001101100011_1_11_110_011_011_0_x_00;
      patterns[1705] = 32'b0101001101100000_1_xx_110_xxx_011_0_1_01;
      patterns[1706] = 32'b0100001101100000_0_xx_110_011_xxx_1_x_xx;
      patterns[1707] = 32'b0000001110001111_1_xx_xxx_xxx_011_0_x_10;
      patterns[1708] = 32'b1000001101100100_1_00_110_100_011_0_x_00;
      patterns[1709] = 32'b1001001101100100_1_01_110_100_011_0_x_00;
      patterns[1710] = 32'b1010001101100100_1_10_110_100_011_0_x_00;
      patterns[1711] = 32'b1011001101100100_1_11_110_100_011_0_x_00;
      patterns[1712] = 32'b0101001101100000_1_xx_110_xxx_011_0_1_01;
      patterns[1713] = 32'b0100001101100000_0_xx_110_011_xxx_1_x_xx;
      patterns[1714] = 32'b0000001101111000_1_xx_xxx_xxx_011_0_x_10;
      patterns[1715] = 32'b1000001101100101_1_00_110_101_011_0_x_00;
      patterns[1716] = 32'b1001001101100101_1_01_110_101_011_0_x_00;
      patterns[1717] = 32'b1010001101100101_1_10_110_101_011_0_x_00;
      patterns[1718] = 32'b1011001101100101_1_11_110_101_011_0_x_00;
      patterns[1719] = 32'b0101001101100000_1_xx_110_xxx_011_0_1_01;
      patterns[1720] = 32'b0100001101100000_0_xx_110_011_xxx_1_x_xx;
      patterns[1721] = 32'b0000001101000111_1_xx_xxx_xxx_011_0_x_10;
      patterns[1722] = 32'b1000001101100110_1_00_110_110_011_0_x_00;
      patterns[1723] = 32'b1001001101100110_1_01_110_110_011_0_x_00;
      patterns[1724] = 32'b1010001101100110_1_10_110_110_011_0_x_00;
      patterns[1725] = 32'b1011001101100110_1_11_110_110_011_0_x_00;
      patterns[1726] = 32'b0101001101100000_1_xx_110_xxx_011_0_1_01;
      patterns[1727] = 32'b0100001101100000_0_xx_110_011_xxx_1_x_xx;
      patterns[1728] = 32'b0000001110101001_1_xx_xxx_xxx_011_0_x_10;
      patterns[1729] = 32'b1000001101100111_1_00_110_111_011_0_x_00;
      patterns[1730] = 32'b1001001101100111_1_01_110_111_011_0_x_00;
      patterns[1731] = 32'b1010001101100111_1_10_110_111_011_0_x_00;
      patterns[1732] = 32'b1011001101100111_1_11_110_111_011_0_x_00;
      patterns[1733] = 32'b0101001101100000_1_xx_110_xxx_011_0_1_01;
      patterns[1734] = 32'b0100001101100000_0_xx_110_011_xxx_1_x_xx;
      patterns[1735] = 32'b0000001101100011_1_xx_xxx_xxx_011_0_x_10;
      patterns[1736] = 32'b1000001101110000_1_00_111_000_011_0_x_00;
      patterns[1737] = 32'b1001001101110000_1_01_111_000_011_0_x_00;
      patterns[1738] = 32'b1010001101110000_1_10_111_000_011_0_x_00;
      patterns[1739] = 32'b1011001101110000_1_11_111_000_011_0_x_00;
      patterns[1740] = 32'b0101001101110000_1_xx_111_xxx_011_0_1_01;
      patterns[1741] = 32'b0100001101110000_0_xx_111_011_xxx_1_x_xx;
      patterns[1742] = 32'b0000001110010011_1_xx_xxx_xxx_011_0_x_10;
      patterns[1743] = 32'b1000001101110001_1_00_111_001_011_0_x_00;
      patterns[1744] = 32'b1001001101110001_1_01_111_001_011_0_x_00;
      patterns[1745] = 32'b1010001101110001_1_10_111_001_011_0_x_00;
      patterns[1746] = 32'b1011001101110001_1_11_111_001_011_0_x_00;
      patterns[1747] = 32'b0101001101110000_1_xx_111_xxx_011_0_1_01;
      patterns[1748] = 32'b0100001101110000_0_xx_111_011_xxx_1_x_xx;
      patterns[1749] = 32'b0000001110001011_1_xx_xxx_xxx_011_0_x_10;
      patterns[1750] = 32'b1000001101110010_1_00_111_010_011_0_x_00;
      patterns[1751] = 32'b1001001101110010_1_01_111_010_011_0_x_00;
      patterns[1752] = 32'b1010001101110010_1_10_111_010_011_0_x_00;
      patterns[1753] = 32'b1011001101110010_1_11_111_010_011_0_x_00;
      patterns[1754] = 32'b0101001101110000_1_xx_111_xxx_011_0_1_01;
      patterns[1755] = 32'b0100001101110000_0_xx_111_011_xxx_1_x_xx;
      patterns[1756] = 32'b0000001101010000_1_xx_xxx_xxx_011_0_x_10;
      patterns[1757] = 32'b1000001101110011_1_00_111_011_011_0_x_00;
      patterns[1758] = 32'b1001001101110011_1_01_111_011_011_0_x_00;
      patterns[1759] = 32'b1010001101110011_1_10_111_011_011_0_x_00;
      patterns[1760] = 32'b1011001101110011_1_11_111_011_011_0_x_00;
      patterns[1761] = 32'b0101001101110000_1_xx_111_xxx_011_0_1_01;
      patterns[1762] = 32'b0100001101110000_0_xx_111_011_xxx_1_x_xx;
      patterns[1763] = 32'b0000001100100000_1_xx_xxx_xxx_011_0_x_10;
      patterns[1764] = 32'b1000001101110100_1_00_111_100_011_0_x_00;
      patterns[1765] = 32'b1001001101110100_1_01_111_100_011_0_x_00;
      patterns[1766] = 32'b1010001101110100_1_10_111_100_011_0_x_00;
      patterns[1767] = 32'b1011001101110100_1_11_111_100_011_0_x_00;
      patterns[1768] = 32'b0101001101110000_1_xx_111_xxx_011_0_1_01;
      patterns[1769] = 32'b0100001101110000_0_xx_111_011_xxx_1_x_xx;
      patterns[1770] = 32'b0000001101000100_1_xx_xxx_xxx_011_0_x_10;
      patterns[1771] = 32'b1000001101110101_1_00_111_101_011_0_x_00;
      patterns[1772] = 32'b1001001101110101_1_01_111_101_011_0_x_00;
      patterns[1773] = 32'b1010001101110101_1_10_111_101_011_0_x_00;
      patterns[1774] = 32'b1011001101110101_1_11_111_101_011_0_x_00;
      patterns[1775] = 32'b0101001101110000_1_xx_111_xxx_011_0_1_01;
      patterns[1776] = 32'b0100001101110000_0_xx_111_011_xxx_1_x_xx;
      patterns[1777] = 32'b0000001110100011_1_xx_xxx_xxx_011_0_x_10;
      patterns[1778] = 32'b1000001101110110_1_00_111_110_011_0_x_00;
      patterns[1779] = 32'b1001001101110110_1_01_111_110_011_0_x_00;
      patterns[1780] = 32'b1010001101110110_1_10_111_110_011_0_x_00;
      patterns[1781] = 32'b1011001101110110_1_11_111_110_011_0_x_00;
      patterns[1782] = 32'b0101001101110000_1_xx_111_xxx_011_0_1_01;
      patterns[1783] = 32'b0100001101110000_0_xx_111_011_xxx_1_x_xx;
      patterns[1784] = 32'b0000001101011101_1_xx_xxx_xxx_011_0_x_10;
      patterns[1785] = 32'b1000001101110111_1_00_111_111_011_0_x_00;
      patterns[1786] = 32'b1001001101110111_1_01_111_111_011_0_x_00;
      patterns[1787] = 32'b1010001101110111_1_10_111_111_011_0_x_00;
      patterns[1788] = 32'b1011001101110111_1_11_111_111_011_0_x_00;
      patterns[1789] = 32'b0101001101110000_1_xx_111_xxx_011_0_1_01;
      patterns[1790] = 32'b0100001101110000_0_xx_111_011_xxx_1_x_xx;
      patterns[1791] = 32'b0000001111000010_1_xx_xxx_xxx_011_0_x_10;
      patterns[1792] = 32'b1000010000000000_1_00_000_000_100_0_x_00;
      patterns[1793] = 32'b1001010000000000_1_01_000_000_100_0_x_00;
      patterns[1794] = 32'b1010010000000000_1_10_000_000_100_0_x_00;
      patterns[1795] = 32'b1011010000000000_1_11_000_000_100_0_x_00;
      patterns[1796] = 32'b0101010000000000_1_xx_000_xxx_100_0_1_01;
      patterns[1797] = 32'b0100010000000000_0_xx_000_100_xxx_1_x_xx;
      patterns[1798] = 32'b0000010011001110_1_xx_xxx_xxx_100_0_x_10;
      patterns[1799] = 32'b1000010000000001_1_00_000_001_100_0_x_00;
      patterns[1800] = 32'b1001010000000001_1_01_000_001_100_0_x_00;
      patterns[1801] = 32'b1010010000000001_1_10_000_001_100_0_x_00;
      patterns[1802] = 32'b1011010000000001_1_11_000_001_100_0_x_00;
      patterns[1803] = 32'b0101010000000000_1_xx_000_xxx_100_0_1_01;
      patterns[1804] = 32'b0100010000000000_0_xx_000_100_xxx_1_x_xx;
      patterns[1805] = 32'b0000010011111110_1_xx_xxx_xxx_100_0_x_10;
      patterns[1806] = 32'b1000010000000010_1_00_000_010_100_0_x_00;
      patterns[1807] = 32'b1001010000000010_1_01_000_010_100_0_x_00;
      patterns[1808] = 32'b1010010000000010_1_10_000_010_100_0_x_00;
      patterns[1809] = 32'b1011010000000010_1_11_000_010_100_0_x_00;
      patterns[1810] = 32'b0101010000000000_1_xx_000_xxx_100_0_1_01;
      patterns[1811] = 32'b0100010000000000_0_xx_000_100_xxx_1_x_xx;
      patterns[1812] = 32'b0000010000101111_1_xx_xxx_xxx_100_0_x_10;
      patterns[1813] = 32'b1000010000000011_1_00_000_011_100_0_x_00;
      patterns[1814] = 32'b1001010000000011_1_01_000_011_100_0_x_00;
      patterns[1815] = 32'b1010010000000011_1_10_000_011_100_0_x_00;
      patterns[1816] = 32'b1011010000000011_1_11_000_011_100_0_x_00;
      patterns[1817] = 32'b0101010000000000_1_xx_000_xxx_100_0_1_01;
      patterns[1818] = 32'b0100010000000000_0_xx_000_100_xxx_1_x_xx;
      patterns[1819] = 32'b0000010010001111_1_xx_xxx_xxx_100_0_x_10;
      patterns[1820] = 32'b1000010000000100_1_00_000_100_100_0_x_00;
      patterns[1821] = 32'b1001010000000100_1_01_000_100_100_0_x_00;
      patterns[1822] = 32'b1010010000000100_1_10_000_100_100_0_x_00;
      patterns[1823] = 32'b1011010000000100_1_11_000_100_100_0_x_00;
      patterns[1824] = 32'b0101010000000000_1_xx_000_xxx_100_0_1_01;
      patterns[1825] = 32'b0100010000000000_0_xx_000_100_xxx_1_x_xx;
      patterns[1826] = 32'b0000010000011001_1_xx_xxx_xxx_100_0_x_10;
      patterns[1827] = 32'b1000010000000101_1_00_000_101_100_0_x_00;
      patterns[1828] = 32'b1001010000000101_1_01_000_101_100_0_x_00;
      patterns[1829] = 32'b1010010000000101_1_10_000_101_100_0_x_00;
      patterns[1830] = 32'b1011010000000101_1_11_000_101_100_0_x_00;
      patterns[1831] = 32'b0101010000000000_1_xx_000_xxx_100_0_1_01;
      patterns[1832] = 32'b0100010000000000_0_xx_000_100_xxx_1_x_xx;
      patterns[1833] = 32'b0000010010001000_1_xx_xxx_xxx_100_0_x_10;
      patterns[1834] = 32'b1000010000000110_1_00_000_110_100_0_x_00;
      patterns[1835] = 32'b1001010000000110_1_01_000_110_100_0_x_00;
      patterns[1836] = 32'b1010010000000110_1_10_000_110_100_0_x_00;
      patterns[1837] = 32'b1011010000000110_1_11_000_110_100_0_x_00;
      patterns[1838] = 32'b0101010000000000_1_xx_000_xxx_100_0_1_01;
      patterns[1839] = 32'b0100010000000000_0_xx_000_100_xxx_1_x_xx;
      patterns[1840] = 32'b0000010010110010_1_xx_xxx_xxx_100_0_x_10;
      patterns[1841] = 32'b1000010000000111_1_00_000_111_100_0_x_00;
      patterns[1842] = 32'b1001010000000111_1_01_000_111_100_0_x_00;
      patterns[1843] = 32'b1010010000000111_1_10_000_111_100_0_x_00;
      patterns[1844] = 32'b1011010000000111_1_11_000_111_100_0_x_00;
      patterns[1845] = 32'b0101010000000000_1_xx_000_xxx_100_0_1_01;
      patterns[1846] = 32'b0100010000000000_0_xx_000_100_xxx_1_x_xx;
      patterns[1847] = 32'b0000010000101110_1_xx_xxx_xxx_100_0_x_10;
      patterns[1848] = 32'b1000010000010000_1_00_001_000_100_0_x_00;
      patterns[1849] = 32'b1001010000010000_1_01_001_000_100_0_x_00;
      patterns[1850] = 32'b1010010000010000_1_10_001_000_100_0_x_00;
      patterns[1851] = 32'b1011010000010000_1_11_001_000_100_0_x_00;
      patterns[1852] = 32'b0101010000010000_1_xx_001_xxx_100_0_1_01;
      patterns[1853] = 32'b0100010000010000_0_xx_001_100_xxx_1_x_xx;
      patterns[1854] = 32'b0000010011111110_1_xx_xxx_xxx_100_0_x_10;
      patterns[1855] = 32'b1000010000010001_1_00_001_001_100_0_x_00;
      patterns[1856] = 32'b1001010000010001_1_01_001_001_100_0_x_00;
      patterns[1857] = 32'b1010010000010001_1_10_001_001_100_0_x_00;
      patterns[1858] = 32'b1011010000010001_1_11_001_001_100_0_x_00;
      patterns[1859] = 32'b0101010000010000_1_xx_001_xxx_100_0_1_01;
      patterns[1860] = 32'b0100010000010000_0_xx_001_100_xxx_1_x_xx;
      patterns[1861] = 32'b0000010011101010_1_xx_xxx_xxx_100_0_x_10;
      patterns[1862] = 32'b1000010000010010_1_00_001_010_100_0_x_00;
      patterns[1863] = 32'b1001010000010010_1_01_001_010_100_0_x_00;
      patterns[1864] = 32'b1010010000010010_1_10_001_010_100_0_x_00;
      patterns[1865] = 32'b1011010000010010_1_11_001_010_100_0_x_00;
      patterns[1866] = 32'b0101010000010000_1_xx_001_xxx_100_0_1_01;
      patterns[1867] = 32'b0100010000010000_0_xx_001_100_xxx_1_x_xx;
      patterns[1868] = 32'b0000010000110000_1_xx_xxx_xxx_100_0_x_10;
      patterns[1869] = 32'b1000010000010011_1_00_001_011_100_0_x_00;
      patterns[1870] = 32'b1001010000010011_1_01_001_011_100_0_x_00;
      patterns[1871] = 32'b1010010000010011_1_10_001_011_100_0_x_00;
      patterns[1872] = 32'b1011010000010011_1_11_001_011_100_0_x_00;
      patterns[1873] = 32'b0101010000010000_1_xx_001_xxx_100_0_1_01;
      patterns[1874] = 32'b0100010000010000_0_xx_001_100_xxx_1_x_xx;
      patterns[1875] = 32'b0000010001100111_1_xx_xxx_xxx_100_0_x_10;
      patterns[1876] = 32'b1000010000010100_1_00_001_100_100_0_x_00;
      patterns[1877] = 32'b1001010000010100_1_01_001_100_100_0_x_00;
      patterns[1878] = 32'b1010010000010100_1_10_001_100_100_0_x_00;
      patterns[1879] = 32'b1011010000010100_1_11_001_100_100_0_x_00;
      patterns[1880] = 32'b0101010000010000_1_xx_001_xxx_100_0_1_01;
      patterns[1881] = 32'b0100010000010000_0_xx_001_100_xxx_1_x_xx;
      patterns[1882] = 32'b0000010001011101_1_xx_xxx_xxx_100_0_x_10;
      patterns[1883] = 32'b1000010000010101_1_00_001_101_100_0_x_00;
      patterns[1884] = 32'b1001010000010101_1_01_001_101_100_0_x_00;
      patterns[1885] = 32'b1010010000010101_1_10_001_101_100_0_x_00;
      patterns[1886] = 32'b1011010000010101_1_11_001_101_100_0_x_00;
      patterns[1887] = 32'b0101010000010000_1_xx_001_xxx_100_0_1_01;
      patterns[1888] = 32'b0100010000010000_0_xx_001_100_xxx_1_x_xx;
      patterns[1889] = 32'b0000010001011011_1_xx_xxx_xxx_100_0_x_10;
      patterns[1890] = 32'b1000010000010110_1_00_001_110_100_0_x_00;
      patterns[1891] = 32'b1001010000010110_1_01_001_110_100_0_x_00;
      patterns[1892] = 32'b1010010000010110_1_10_001_110_100_0_x_00;
      patterns[1893] = 32'b1011010000010110_1_11_001_110_100_0_x_00;
      patterns[1894] = 32'b0101010000010000_1_xx_001_xxx_100_0_1_01;
      patterns[1895] = 32'b0100010000010000_0_xx_001_100_xxx_1_x_xx;
      patterns[1896] = 32'b0000010010011101_1_xx_xxx_xxx_100_0_x_10;
      patterns[1897] = 32'b1000010000010111_1_00_001_111_100_0_x_00;
      patterns[1898] = 32'b1001010000010111_1_01_001_111_100_0_x_00;
      patterns[1899] = 32'b1010010000010111_1_10_001_111_100_0_x_00;
      patterns[1900] = 32'b1011010000010111_1_11_001_111_100_0_x_00;
      patterns[1901] = 32'b0101010000010000_1_xx_001_xxx_100_0_1_01;
      patterns[1902] = 32'b0100010000010000_0_xx_001_100_xxx_1_x_xx;
      patterns[1903] = 32'b0000010001011011_1_xx_xxx_xxx_100_0_x_10;
      patterns[1904] = 32'b1000010000100000_1_00_010_000_100_0_x_00;
      patterns[1905] = 32'b1001010000100000_1_01_010_000_100_0_x_00;
      patterns[1906] = 32'b1010010000100000_1_10_010_000_100_0_x_00;
      patterns[1907] = 32'b1011010000100000_1_11_010_000_100_0_x_00;
      patterns[1908] = 32'b0101010000100000_1_xx_010_xxx_100_0_1_01;
      patterns[1909] = 32'b0100010000100000_0_xx_010_100_xxx_1_x_xx;
      patterns[1910] = 32'b0000010010110101_1_xx_xxx_xxx_100_0_x_10;
      patterns[1911] = 32'b1000010000100001_1_00_010_001_100_0_x_00;
      patterns[1912] = 32'b1001010000100001_1_01_010_001_100_0_x_00;
      patterns[1913] = 32'b1010010000100001_1_10_010_001_100_0_x_00;
      patterns[1914] = 32'b1011010000100001_1_11_010_001_100_0_x_00;
      patterns[1915] = 32'b0101010000100000_1_xx_010_xxx_100_0_1_01;
      patterns[1916] = 32'b0100010000100000_0_xx_010_100_xxx_1_x_xx;
      patterns[1917] = 32'b0000010001100000_1_xx_xxx_xxx_100_0_x_10;
      patterns[1918] = 32'b1000010000100010_1_00_010_010_100_0_x_00;
      patterns[1919] = 32'b1001010000100010_1_01_010_010_100_0_x_00;
      patterns[1920] = 32'b1010010000100010_1_10_010_010_100_0_x_00;
      patterns[1921] = 32'b1011010000100010_1_11_010_010_100_0_x_00;
      patterns[1922] = 32'b0101010000100000_1_xx_010_xxx_100_0_1_01;
      patterns[1923] = 32'b0100010000100000_0_xx_010_100_xxx_1_x_xx;
      patterns[1924] = 32'b0000010000111100_1_xx_xxx_xxx_100_0_x_10;
      patterns[1925] = 32'b1000010000100011_1_00_010_011_100_0_x_00;
      patterns[1926] = 32'b1001010000100011_1_01_010_011_100_0_x_00;
      patterns[1927] = 32'b1010010000100011_1_10_010_011_100_0_x_00;
      patterns[1928] = 32'b1011010000100011_1_11_010_011_100_0_x_00;
      patterns[1929] = 32'b0101010000100000_1_xx_010_xxx_100_0_1_01;
      patterns[1930] = 32'b0100010000100000_0_xx_010_100_xxx_1_x_xx;
      patterns[1931] = 32'b0000010001110101_1_xx_xxx_xxx_100_0_x_10;
      patterns[1932] = 32'b1000010000100100_1_00_010_100_100_0_x_00;
      patterns[1933] = 32'b1001010000100100_1_01_010_100_100_0_x_00;
      patterns[1934] = 32'b1010010000100100_1_10_010_100_100_0_x_00;
      patterns[1935] = 32'b1011010000100100_1_11_010_100_100_0_x_00;
      patterns[1936] = 32'b0101010000100000_1_xx_010_xxx_100_0_1_01;
      patterns[1937] = 32'b0100010000100000_0_xx_010_100_xxx_1_x_xx;
      patterns[1938] = 32'b0000010011100110_1_xx_xxx_xxx_100_0_x_10;
      patterns[1939] = 32'b1000010000100101_1_00_010_101_100_0_x_00;
      patterns[1940] = 32'b1001010000100101_1_01_010_101_100_0_x_00;
      patterns[1941] = 32'b1010010000100101_1_10_010_101_100_0_x_00;
      patterns[1942] = 32'b1011010000100101_1_11_010_101_100_0_x_00;
      patterns[1943] = 32'b0101010000100000_1_xx_010_xxx_100_0_1_01;
      patterns[1944] = 32'b0100010000100000_0_xx_010_100_xxx_1_x_xx;
      patterns[1945] = 32'b0000010000111011_1_xx_xxx_xxx_100_0_x_10;
      patterns[1946] = 32'b1000010000100110_1_00_010_110_100_0_x_00;
      patterns[1947] = 32'b1001010000100110_1_01_010_110_100_0_x_00;
      patterns[1948] = 32'b1010010000100110_1_10_010_110_100_0_x_00;
      patterns[1949] = 32'b1011010000100110_1_11_010_110_100_0_x_00;
      patterns[1950] = 32'b0101010000100000_1_xx_010_xxx_100_0_1_01;
      patterns[1951] = 32'b0100010000100000_0_xx_010_100_xxx_1_x_xx;
      patterns[1952] = 32'b0000010000110111_1_xx_xxx_xxx_100_0_x_10;
      patterns[1953] = 32'b1000010000100111_1_00_010_111_100_0_x_00;
      patterns[1954] = 32'b1001010000100111_1_01_010_111_100_0_x_00;
      patterns[1955] = 32'b1010010000100111_1_10_010_111_100_0_x_00;
      patterns[1956] = 32'b1011010000100111_1_11_010_111_100_0_x_00;
      patterns[1957] = 32'b0101010000100000_1_xx_010_xxx_100_0_1_01;
      patterns[1958] = 32'b0100010000100000_0_xx_010_100_xxx_1_x_xx;
      patterns[1959] = 32'b0000010001111011_1_xx_xxx_xxx_100_0_x_10;
      patterns[1960] = 32'b1000010000110000_1_00_011_000_100_0_x_00;
      patterns[1961] = 32'b1001010000110000_1_01_011_000_100_0_x_00;
      patterns[1962] = 32'b1010010000110000_1_10_011_000_100_0_x_00;
      patterns[1963] = 32'b1011010000110000_1_11_011_000_100_0_x_00;
      patterns[1964] = 32'b0101010000110000_1_xx_011_xxx_100_0_1_01;
      patterns[1965] = 32'b0100010000110000_0_xx_011_100_xxx_1_x_xx;
      patterns[1966] = 32'b0000010010011000_1_xx_xxx_xxx_100_0_x_10;
      patterns[1967] = 32'b1000010000110001_1_00_011_001_100_0_x_00;
      patterns[1968] = 32'b1001010000110001_1_01_011_001_100_0_x_00;
      patterns[1969] = 32'b1010010000110001_1_10_011_001_100_0_x_00;
      patterns[1970] = 32'b1011010000110001_1_11_011_001_100_0_x_00;
      patterns[1971] = 32'b0101010000110000_1_xx_011_xxx_100_0_1_01;
      patterns[1972] = 32'b0100010000110000_0_xx_011_100_xxx_1_x_xx;
      patterns[1973] = 32'b0000010000110000_1_xx_xxx_xxx_100_0_x_10;
      patterns[1974] = 32'b1000010000110010_1_00_011_010_100_0_x_00;
      patterns[1975] = 32'b1001010000110010_1_01_011_010_100_0_x_00;
      patterns[1976] = 32'b1010010000110010_1_10_011_010_100_0_x_00;
      patterns[1977] = 32'b1011010000110010_1_11_011_010_100_0_x_00;
      patterns[1978] = 32'b0101010000110000_1_xx_011_xxx_100_0_1_01;
      patterns[1979] = 32'b0100010000110000_0_xx_011_100_xxx_1_x_xx;
      patterns[1980] = 32'b0000010000111100_1_xx_xxx_xxx_100_0_x_10;
      patterns[1981] = 32'b1000010000110011_1_00_011_011_100_0_x_00;
      patterns[1982] = 32'b1001010000110011_1_01_011_011_100_0_x_00;
      patterns[1983] = 32'b1010010000110011_1_10_011_011_100_0_x_00;
      patterns[1984] = 32'b1011010000110011_1_11_011_011_100_0_x_00;
      patterns[1985] = 32'b0101010000110000_1_xx_011_xxx_100_0_1_01;
      patterns[1986] = 32'b0100010000110000_0_xx_011_100_xxx_1_x_xx;
      patterns[1987] = 32'b0000010001011010_1_xx_xxx_xxx_100_0_x_10;
      patterns[1988] = 32'b1000010000110100_1_00_011_100_100_0_x_00;
      patterns[1989] = 32'b1001010000110100_1_01_011_100_100_0_x_00;
      patterns[1990] = 32'b1010010000110100_1_10_011_100_100_0_x_00;
      patterns[1991] = 32'b1011010000110100_1_11_011_100_100_0_x_00;
      patterns[1992] = 32'b0101010000110000_1_xx_011_xxx_100_0_1_01;
      patterns[1993] = 32'b0100010000110000_0_xx_011_100_xxx_1_x_xx;
      patterns[1994] = 32'b0000010000010110_1_xx_xxx_xxx_100_0_x_10;
      patterns[1995] = 32'b1000010000110101_1_00_011_101_100_0_x_00;
      patterns[1996] = 32'b1001010000110101_1_01_011_101_100_0_x_00;
      patterns[1997] = 32'b1010010000110101_1_10_011_101_100_0_x_00;
      patterns[1998] = 32'b1011010000110101_1_11_011_101_100_0_x_00;
      patterns[1999] = 32'b0101010000110000_1_xx_011_xxx_100_0_1_01;
      patterns[2000] = 32'b0100010000110000_0_xx_011_100_xxx_1_x_xx;
      patterns[2001] = 32'b0000010011000110_1_xx_xxx_xxx_100_0_x_10;
      patterns[2002] = 32'b1000010000110110_1_00_011_110_100_0_x_00;
      patterns[2003] = 32'b1001010000110110_1_01_011_110_100_0_x_00;
      patterns[2004] = 32'b1010010000110110_1_10_011_110_100_0_x_00;
      patterns[2005] = 32'b1011010000110110_1_11_011_110_100_0_x_00;
      patterns[2006] = 32'b0101010000110000_1_xx_011_xxx_100_0_1_01;
      patterns[2007] = 32'b0100010000110000_0_xx_011_100_xxx_1_x_xx;
      patterns[2008] = 32'b0000010000111110_1_xx_xxx_xxx_100_0_x_10;
      patterns[2009] = 32'b1000010000110111_1_00_011_111_100_0_x_00;
      patterns[2010] = 32'b1001010000110111_1_01_011_111_100_0_x_00;
      patterns[2011] = 32'b1010010000110111_1_10_011_111_100_0_x_00;
      patterns[2012] = 32'b1011010000110111_1_11_011_111_100_0_x_00;
      patterns[2013] = 32'b0101010000110000_1_xx_011_xxx_100_0_1_01;
      patterns[2014] = 32'b0100010000110000_0_xx_011_100_xxx_1_x_xx;
      patterns[2015] = 32'b0000010000110111_1_xx_xxx_xxx_100_0_x_10;
      patterns[2016] = 32'b1000010001000000_1_00_100_000_100_0_x_00;
      patterns[2017] = 32'b1001010001000000_1_01_100_000_100_0_x_00;
      patterns[2018] = 32'b1010010001000000_1_10_100_000_100_0_x_00;
      patterns[2019] = 32'b1011010001000000_1_11_100_000_100_0_x_00;
      patterns[2020] = 32'b0101010001000000_1_xx_100_xxx_100_0_1_01;
      patterns[2021] = 32'b0100010001000000_0_xx_100_100_xxx_1_x_xx;
      patterns[2022] = 32'b0000010010000110_1_xx_xxx_xxx_100_0_x_10;
      patterns[2023] = 32'b1000010001000001_1_00_100_001_100_0_x_00;
      patterns[2024] = 32'b1001010001000001_1_01_100_001_100_0_x_00;
      patterns[2025] = 32'b1010010001000001_1_10_100_001_100_0_x_00;
      patterns[2026] = 32'b1011010001000001_1_11_100_001_100_0_x_00;
      patterns[2027] = 32'b0101010001000000_1_xx_100_xxx_100_0_1_01;
      patterns[2028] = 32'b0100010001000000_0_xx_100_100_xxx_1_x_xx;
      patterns[2029] = 32'b0000010010000100_1_xx_xxx_xxx_100_0_x_10;
      patterns[2030] = 32'b1000010001000010_1_00_100_010_100_0_x_00;
      patterns[2031] = 32'b1001010001000010_1_01_100_010_100_0_x_00;
      patterns[2032] = 32'b1010010001000010_1_10_100_010_100_0_x_00;
      patterns[2033] = 32'b1011010001000010_1_11_100_010_100_0_x_00;
      patterns[2034] = 32'b0101010001000000_1_xx_100_xxx_100_0_1_01;
      patterns[2035] = 32'b0100010001000000_0_xx_100_100_xxx_1_x_xx;
      patterns[2036] = 32'b0000010001010010_1_xx_xxx_xxx_100_0_x_10;
      patterns[2037] = 32'b1000010001000011_1_00_100_011_100_0_x_00;
      patterns[2038] = 32'b1001010001000011_1_01_100_011_100_0_x_00;
      patterns[2039] = 32'b1010010001000011_1_10_100_011_100_0_x_00;
      patterns[2040] = 32'b1011010001000011_1_11_100_011_100_0_x_00;
      patterns[2041] = 32'b0101010001000000_1_xx_100_xxx_100_0_1_01;
      patterns[2042] = 32'b0100010001000000_0_xx_100_100_xxx_1_x_xx;
      patterns[2043] = 32'b0000010001001111_1_xx_xxx_xxx_100_0_x_10;
      patterns[2044] = 32'b1000010001000100_1_00_100_100_100_0_x_00;
      patterns[2045] = 32'b1001010001000100_1_01_100_100_100_0_x_00;
      patterns[2046] = 32'b1010010001000100_1_10_100_100_100_0_x_00;
      patterns[2047] = 32'b1011010001000100_1_11_100_100_100_0_x_00;
      patterns[2048] = 32'b0101010001000000_1_xx_100_xxx_100_0_1_01;
      patterns[2049] = 32'b0100010001000000_0_xx_100_100_xxx_1_x_xx;
      patterns[2050] = 32'b0000010000001001_1_xx_xxx_xxx_100_0_x_10;
      patterns[2051] = 32'b1000010001000101_1_00_100_101_100_0_x_00;
      patterns[2052] = 32'b1001010001000101_1_01_100_101_100_0_x_00;
      patterns[2053] = 32'b1010010001000101_1_10_100_101_100_0_x_00;
      patterns[2054] = 32'b1011010001000101_1_11_100_101_100_0_x_00;
      patterns[2055] = 32'b0101010001000000_1_xx_100_xxx_100_0_1_01;
      patterns[2056] = 32'b0100010001000000_0_xx_100_100_xxx_1_x_xx;
      patterns[2057] = 32'b0000010010000010_1_xx_xxx_xxx_100_0_x_10;
      patterns[2058] = 32'b1000010001000110_1_00_100_110_100_0_x_00;
      patterns[2059] = 32'b1001010001000110_1_01_100_110_100_0_x_00;
      patterns[2060] = 32'b1010010001000110_1_10_100_110_100_0_x_00;
      patterns[2061] = 32'b1011010001000110_1_11_100_110_100_0_x_00;
      patterns[2062] = 32'b0101010001000000_1_xx_100_xxx_100_0_1_01;
      patterns[2063] = 32'b0100010001000000_0_xx_100_100_xxx_1_x_xx;
      patterns[2064] = 32'b0000010011011101_1_xx_xxx_xxx_100_0_x_10;
      patterns[2065] = 32'b1000010001000111_1_00_100_111_100_0_x_00;
      patterns[2066] = 32'b1001010001000111_1_01_100_111_100_0_x_00;
      patterns[2067] = 32'b1010010001000111_1_10_100_111_100_0_x_00;
      patterns[2068] = 32'b1011010001000111_1_11_100_111_100_0_x_00;
      patterns[2069] = 32'b0101010001000000_1_xx_100_xxx_100_0_1_01;
      patterns[2070] = 32'b0100010001000000_0_xx_100_100_xxx_1_x_xx;
      patterns[2071] = 32'b0000010000011100_1_xx_xxx_xxx_100_0_x_10;
      patterns[2072] = 32'b1000010001010000_1_00_101_000_100_0_x_00;
      patterns[2073] = 32'b1001010001010000_1_01_101_000_100_0_x_00;
      patterns[2074] = 32'b1010010001010000_1_10_101_000_100_0_x_00;
      patterns[2075] = 32'b1011010001010000_1_11_101_000_100_0_x_00;
      patterns[2076] = 32'b0101010001010000_1_xx_101_xxx_100_0_1_01;
      patterns[2077] = 32'b0100010001010000_0_xx_101_100_xxx_1_x_xx;
      patterns[2078] = 32'b0000010010111111_1_xx_xxx_xxx_100_0_x_10;
      patterns[2079] = 32'b1000010001010001_1_00_101_001_100_0_x_00;
      patterns[2080] = 32'b1001010001010001_1_01_101_001_100_0_x_00;
      patterns[2081] = 32'b1010010001010001_1_10_101_001_100_0_x_00;
      patterns[2082] = 32'b1011010001010001_1_11_101_001_100_0_x_00;
      patterns[2083] = 32'b0101010001010000_1_xx_101_xxx_100_0_1_01;
      patterns[2084] = 32'b0100010001010000_0_xx_101_100_xxx_1_x_xx;
      patterns[2085] = 32'b0000010000110100_1_xx_xxx_xxx_100_0_x_10;
      patterns[2086] = 32'b1000010001010010_1_00_101_010_100_0_x_00;
      patterns[2087] = 32'b1001010001010010_1_01_101_010_100_0_x_00;
      patterns[2088] = 32'b1010010001010010_1_10_101_010_100_0_x_00;
      patterns[2089] = 32'b1011010001010010_1_11_101_010_100_0_x_00;
      patterns[2090] = 32'b0101010001010000_1_xx_101_xxx_100_0_1_01;
      patterns[2091] = 32'b0100010001010000_0_xx_101_100_xxx_1_x_xx;
      patterns[2092] = 32'b0000010010000001_1_xx_xxx_xxx_100_0_x_10;
      patterns[2093] = 32'b1000010001010011_1_00_101_011_100_0_x_00;
      patterns[2094] = 32'b1001010001010011_1_01_101_011_100_0_x_00;
      patterns[2095] = 32'b1010010001010011_1_10_101_011_100_0_x_00;
      patterns[2096] = 32'b1011010001010011_1_11_101_011_100_0_x_00;
      patterns[2097] = 32'b0101010001010000_1_xx_101_xxx_100_0_1_01;
      patterns[2098] = 32'b0100010001010000_0_xx_101_100_xxx_1_x_xx;
      patterns[2099] = 32'b0000010011001011_1_xx_xxx_xxx_100_0_x_10;
      patterns[2100] = 32'b1000010001010100_1_00_101_100_100_0_x_00;
      patterns[2101] = 32'b1001010001010100_1_01_101_100_100_0_x_00;
      patterns[2102] = 32'b1010010001010100_1_10_101_100_100_0_x_00;
      patterns[2103] = 32'b1011010001010100_1_11_101_100_100_0_x_00;
      patterns[2104] = 32'b0101010001010000_1_xx_101_xxx_100_0_1_01;
      patterns[2105] = 32'b0100010001010000_0_xx_101_100_xxx_1_x_xx;
      patterns[2106] = 32'b0000010010001101_1_xx_xxx_xxx_100_0_x_10;
      patterns[2107] = 32'b1000010001010101_1_00_101_101_100_0_x_00;
      patterns[2108] = 32'b1001010001010101_1_01_101_101_100_0_x_00;
      patterns[2109] = 32'b1010010001010101_1_10_101_101_100_0_x_00;
      patterns[2110] = 32'b1011010001010101_1_11_101_101_100_0_x_00;
      patterns[2111] = 32'b0101010001010000_1_xx_101_xxx_100_0_1_01;
      patterns[2112] = 32'b0100010001010000_0_xx_101_100_xxx_1_x_xx;
      patterns[2113] = 32'b0000010010000010_1_xx_xxx_xxx_100_0_x_10;
      patterns[2114] = 32'b1000010001010110_1_00_101_110_100_0_x_00;
      patterns[2115] = 32'b1001010001010110_1_01_101_110_100_0_x_00;
      patterns[2116] = 32'b1010010001010110_1_10_101_110_100_0_x_00;
      patterns[2117] = 32'b1011010001010110_1_11_101_110_100_0_x_00;
      patterns[2118] = 32'b0101010001010000_1_xx_101_xxx_100_0_1_01;
      patterns[2119] = 32'b0100010001010000_0_xx_101_100_xxx_1_x_xx;
      patterns[2120] = 32'b0000010011010011_1_xx_xxx_xxx_100_0_x_10;
      patterns[2121] = 32'b1000010001010111_1_00_101_111_100_0_x_00;
      patterns[2122] = 32'b1001010001010111_1_01_101_111_100_0_x_00;
      patterns[2123] = 32'b1010010001010111_1_10_101_111_100_0_x_00;
      patterns[2124] = 32'b1011010001010111_1_11_101_111_100_0_x_00;
      patterns[2125] = 32'b0101010001010000_1_xx_101_xxx_100_0_1_01;
      patterns[2126] = 32'b0100010001010000_0_xx_101_100_xxx_1_x_xx;
      patterns[2127] = 32'b0000010011011101_1_xx_xxx_xxx_100_0_x_10;
      patterns[2128] = 32'b1000010001100000_1_00_110_000_100_0_x_00;
      patterns[2129] = 32'b1001010001100000_1_01_110_000_100_0_x_00;
      patterns[2130] = 32'b1010010001100000_1_10_110_000_100_0_x_00;
      patterns[2131] = 32'b1011010001100000_1_11_110_000_100_0_x_00;
      patterns[2132] = 32'b0101010001100000_1_xx_110_xxx_100_0_1_01;
      patterns[2133] = 32'b0100010001100000_0_xx_110_100_xxx_1_x_xx;
      patterns[2134] = 32'b0000010001011110_1_xx_xxx_xxx_100_0_x_10;
      patterns[2135] = 32'b1000010001100001_1_00_110_001_100_0_x_00;
      patterns[2136] = 32'b1001010001100001_1_01_110_001_100_0_x_00;
      patterns[2137] = 32'b1010010001100001_1_10_110_001_100_0_x_00;
      patterns[2138] = 32'b1011010001100001_1_11_110_001_100_0_x_00;
      patterns[2139] = 32'b0101010001100000_1_xx_110_xxx_100_0_1_01;
      patterns[2140] = 32'b0100010001100000_0_xx_110_100_xxx_1_x_xx;
      patterns[2141] = 32'b0000010000111001_1_xx_xxx_xxx_100_0_x_10;
      patterns[2142] = 32'b1000010001100010_1_00_110_010_100_0_x_00;
      patterns[2143] = 32'b1001010001100010_1_01_110_010_100_0_x_00;
      patterns[2144] = 32'b1010010001100010_1_10_110_010_100_0_x_00;
      patterns[2145] = 32'b1011010001100010_1_11_110_010_100_0_x_00;
      patterns[2146] = 32'b0101010001100000_1_xx_110_xxx_100_0_1_01;
      patterns[2147] = 32'b0100010001100000_0_xx_110_100_xxx_1_x_xx;
      patterns[2148] = 32'b0000010001001110_1_xx_xxx_xxx_100_0_x_10;
      patterns[2149] = 32'b1000010001100011_1_00_110_011_100_0_x_00;
      patterns[2150] = 32'b1001010001100011_1_01_110_011_100_0_x_00;
      patterns[2151] = 32'b1010010001100011_1_10_110_011_100_0_x_00;
      patterns[2152] = 32'b1011010001100011_1_11_110_011_100_0_x_00;
      patterns[2153] = 32'b0101010001100000_1_xx_110_xxx_100_0_1_01;
      patterns[2154] = 32'b0100010001100000_0_xx_110_100_xxx_1_x_xx;
      patterns[2155] = 32'b0000010001010011_1_xx_xxx_xxx_100_0_x_10;
      patterns[2156] = 32'b1000010001100100_1_00_110_100_100_0_x_00;
      patterns[2157] = 32'b1001010001100100_1_01_110_100_100_0_x_00;
      patterns[2158] = 32'b1010010001100100_1_10_110_100_100_0_x_00;
      patterns[2159] = 32'b1011010001100100_1_11_110_100_100_0_x_00;
      patterns[2160] = 32'b0101010001100000_1_xx_110_xxx_100_0_1_01;
      patterns[2161] = 32'b0100010001100000_0_xx_110_100_xxx_1_x_xx;
      patterns[2162] = 32'b0000010010110111_1_xx_xxx_xxx_100_0_x_10;
      patterns[2163] = 32'b1000010001100101_1_00_110_101_100_0_x_00;
      patterns[2164] = 32'b1001010001100101_1_01_110_101_100_0_x_00;
      patterns[2165] = 32'b1010010001100101_1_10_110_101_100_0_x_00;
      patterns[2166] = 32'b1011010001100101_1_11_110_101_100_0_x_00;
      patterns[2167] = 32'b0101010001100000_1_xx_110_xxx_100_0_1_01;
      patterns[2168] = 32'b0100010001100000_0_xx_110_100_xxx_1_x_xx;
      patterns[2169] = 32'b0000010000111011_1_xx_xxx_xxx_100_0_x_10;
      patterns[2170] = 32'b1000010001100110_1_00_110_110_100_0_x_00;
      patterns[2171] = 32'b1001010001100110_1_01_110_110_100_0_x_00;
      patterns[2172] = 32'b1010010001100110_1_10_110_110_100_0_x_00;
      patterns[2173] = 32'b1011010001100110_1_11_110_110_100_0_x_00;
      patterns[2174] = 32'b0101010001100000_1_xx_110_xxx_100_0_1_01;
      patterns[2175] = 32'b0100010001100000_0_xx_110_100_xxx_1_x_xx;
      patterns[2176] = 32'b0000010000000111_1_xx_xxx_xxx_100_0_x_10;
      patterns[2177] = 32'b1000010001100111_1_00_110_111_100_0_x_00;
      patterns[2178] = 32'b1001010001100111_1_01_110_111_100_0_x_00;
      patterns[2179] = 32'b1010010001100111_1_10_110_111_100_0_x_00;
      patterns[2180] = 32'b1011010001100111_1_11_110_111_100_0_x_00;
      patterns[2181] = 32'b0101010001100000_1_xx_110_xxx_100_0_1_01;
      patterns[2182] = 32'b0100010001100000_0_xx_110_100_xxx_1_x_xx;
      patterns[2183] = 32'b0000010000110101_1_xx_xxx_xxx_100_0_x_10;
      patterns[2184] = 32'b1000010001110000_1_00_111_000_100_0_x_00;
      patterns[2185] = 32'b1001010001110000_1_01_111_000_100_0_x_00;
      patterns[2186] = 32'b1010010001110000_1_10_111_000_100_0_x_00;
      patterns[2187] = 32'b1011010001110000_1_11_111_000_100_0_x_00;
      patterns[2188] = 32'b0101010001110000_1_xx_111_xxx_100_0_1_01;
      patterns[2189] = 32'b0100010001110000_0_xx_111_100_xxx_1_x_xx;
      patterns[2190] = 32'b0000010010011100_1_xx_xxx_xxx_100_0_x_10;
      patterns[2191] = 32'b1000010001110001_1_00_111_001_100_0_x_00;
      patterns[2192] = 32'b1001010001110001_1_01_111_001_100_0_x_00;
      patterns[2193] = 32'b1010010001110001_1_10_111_001_100_0_x_00;
      patterns[2194] = 32'b1011010001110001_1_11_111_001_100_0_x_00;
      patterns[2195] = 32'b0101010001110000_1_xx_111_xxx_100_0_1_01;
      patterns[2196] = 32'b0100010001110000_0_xx_111_100_xxx_1_x_xx;
      patterns[2197] = 32'b0000010010110101_1_xx_xxx_xxx_100_0_x_10;
      patterns[2198] = 32'b1000010001110010_1_00_111_010_100_0_x_00;
      patterns[2199] = 32'b1001010001110010_1_01_111_010_100_0_x_00;
      patterns[2200] = 32'b1010010001110010_1_10_111_010_100_0_x_00;
      patterns[2201] = 32'b1011010001110010_1_11_111_010_100_0_x_00;
      patterns[2202] = 32'b0101010001110000_1_xx_111_xxx_100_0_1_01;
      patterns[2203] = 32'b0100010001110000_0_xx_111_100_xxx_1_x_xx;
      patterns[2204] = 32'b0000010000110011_1_xx_xxx_xxx_100_0_x_10;
      patterns[2205] = 32'b1000010001110011_1_00_111_011_100_0_x_00;
      patterns[2206] = 32'b1001010001110011_1_01_111_011_100_0_x_00;
      patterns[2207] = 32'b1010010001110011_1_10_111_011_100_0_x_00;
      patterns[2208] = 32'b1011010001110011_1_11_111_011_100_0_x_00;
      patterns[2209] = 32'b0101010001110000_1_xx_111_xxx_100_0_1_01;
      patterns[2210] = 32'b0100010001110000_0_xx_111_100_xxx_1_x_xx;
      patterns[2211] = 32'b0000010010110100_1_xx_xxx_xxx_100_0_x_10;
      patterns[2212] = 32'b1000010001110100_1_00_111_100_100_0_x_00;
      patterns[2213] = 32'b1001010001110100_1_01_111_100_100_0_x_00;
      patterns[2214] = 32'b1010010001110100_1_10_111_100_100_0_x_00;
      patterns[2215] = 32'b1011010001110100_1_11_111_100_100_0_x_00;
      patterns[2216] = 32'b0101010001110000_1_xx_111_xxx_100_0_1_01;
      patterns[2217] = 32'b0100010001110000_0_xx_111_100_xxx_1_x_xx;
      patterns[2218] = 32'b0000010001001000_1_xx_xxx_xxx_100_0_x_10;
      patterns[2219] = 32'b1000010001110101_1_00_111_101_100_0_x_00;
      patterns[2220] = 32'b1001010001110101_1_01_111_101_100_0_x_00;
      patterns[2221] = 32'b1010010001110101_1_10_111_101_100_0_x_00;
      patterns[2222] = 32'b1011010001110101_1_11_111_101_100_0_x_00;
      patterns[2223] = 32'b0101010001110000_1_xx_111_xxx_100_0_1_01;
      patterns[2224] = 32'b0100010001110000_0_xx_111_100_xxx_1_x_xx;
      patterns[2225] = 32'b0000010010111010_1_xx_xxx_xxx_100_0_x_10;
      patterns[2226] = 32'b1000010001110110_1_00_111_110_100_0_x_00;
      patterns[2227] = 32'b1001010001110110_1_01_111_110_100_0_x_00;
      patterns[2228] = 32'b1010010001110110_1_10_111_110_100_0_x_00;
      patterns[2229] = 32'b1011010001110110_1_11_111_110_100_0_x_00;
      patterns[2230] = 32'b0101010001110000_1_xx_111_xxx_100_0_1_01;
      patterns[2231] = 32'b0100010001110000_0_xx_111_100_xxx_1_x_xx;
      patterns[2232] = 32'b0000010000100000_1_xx_xxx_xxx_100_0_x_10;
      patterns[2233] = 32'b1000010001110111_1_00_111_111_100_0_x_00;
      patterns[2234] = 32'b1001010001110111_1_01_111_111_100_0_x_00;
      patterns[2235] = 32'b1010010001110111_1_10_111_111_100_0_x_00;
      patterns[2236] = 32'b1011010001110111_1_11_111_111_100_0_x_00;
      patterns[2237] = 32'b0101010001110000_1_xx_111_xxx_100_0_1_01;
      patterns[2238] = 32'b0100010001110000_0_xx_111_100_xxx_1_x_xx;
      patterns[2239] = 32'b0000010001100110_1_xx_xxx_xxx_100_0_x_10;
      patterns[2240] = 32'b1000010100000000_1_00_000_000_101_0_x_00;
      patterns[2241] = 32'b1001010100000000_1_01_000_000_101_0_x_00;
      patterns[2242] = 32'b1010010100000000_1_10_000_000_101_0_x_00;
      patterns[2243] = 32'b1011010100000000_1_11_000_000_101_0_x_00;
      patterns[2244] = 32'b0101010100000000_1_xx_000_xxx_101_0_1_01;
      patterns[2245] = 32'b0100010100000000_0_xx_000_101_xxx_1_x_xx;
      patterns[2246] = 32'b0000010110100110_1_xx_xxx_xxx_101_0_x_10;
      patterns[2247] = 32'b1000010100000001_1_00_000_001_101_0_x_00;
      patterns[2248] = 32'b1001010100000001_1_01_000_001_101_0_x_00;
      patterns[2249] = 32'b1010010100000001_1_10_000_001_101_0_x_00;
      patterns[2250] = 32'b1011010100000001_1_11_000_001_101_0_x_00;
      patterns[2251] = 32'b0101010100000000_1_xx_000_xxx_101_0_1_01;
      patterns[2252] = 32'b0100010100000000_0_xx_000_101_xxx_1_x_xx;
      patterns[2253] = 32'b0000010101101010_1_xx_xxx_xxx_101_0_x_10;
      patterns[2254] = 32'b1000010100000010_1_00_000_010_101_0_x_00;
      patterns[2255] = 32'b1001010100000010_1_01_000_010_101_0_x_00;
      patterns[2256] = 32'b1010010100000010_1_10_000_010_101_0_x_00;
      patterns[2257] = 32'b1011010100000010_1_11_000_010_101_0_x_00;
      patterns[2258] = 32'b0101010100000000_1_xx_000_xxx_101_0_1_01;
      patterns[2259] = 32'b0100010100000000_0_xx_000_101_xxx_1_x_xx;
      patterns[2260] = 32'b0000010111111101_1_xx_xxx_xxx_101_0_x_10;
      patterns[2261] = 32'b1000010100000011_1_00_000_011_101_0_x_00;
      patterns[2262] = 32'b1001010100000011_1_01_000_011_101_0_x_00;
      patterns[2263] = 32'b1010010100000011_1_10_000_011_101_0_x_00;
      patterns[2264] = 32'b1011010100000011_1_11_000_011_101_0_x_00;
      patterns[2265] = 32'b0101010100000000_1_xx_000_xxx_101_0_1_01;
      patterns[2266] = 32'b0100010100000000_0_xx_000_101_xxx_1_x_xx;
      patterns[2267] = 32'b0000010101010001_1_xx_xxx_xxx_101_0_x_10;
      patterns[2268] = 32'b1000010100000100_1_00_000_100_101_0_x_00;
      patterns[2269] = 32'b1001010100000100_1_01_000_100_101_0_x_00;
      patterns[2270] = 32'b1010010100000100_1_10_000_100_101_0_x_00;
      patterns[2271] = 32'b1011010100000100_1_11_000_100_101_0_x_00;
      patterns[2272] = 32'b0101010100000000_1_xx_000_xxx_101_0_1_01;
      patterns[2273] = 32'b0100010100000000_0_xx_000_101_xxx_1_x_xx;
      patterns[2274] = 32'b0000010100111100_1_xx_xxx_xxx_101_0_x_10;
      patterns[2275] = 32'b1000010100000101_1_00_000_101_101_0_x_00;
      patterns[2276] = 32'b1001010100000101_1_01_000_101_101_0_x_00;
      patterns[2277] = 32'b1010010100000101_1_10_000_101_101_0_x_00;
      patterns[2278] = 32'b1011010100000101_1_11_000_101_101_0_x_00;
      patterns[2279] = 32'b0101010100000000_1_xx_000_xxx_101_0_1_01;
      patterns[2280] = 32'b0100010100000000_0_xx_000_101_xxx_1_x_xx;
      patterns[2281] = 32'b0000010110011101_1_xx_xxx_xxx_101_0_x_10;
      patterns[2282] = 32'b1000010100000110_1_00_000_110_101_0_x_00;
      patterns[2283] = 32'b1001010100000110_1_01_000_110_101_0_x_00;
      patterns[2284] = 32'b1010010100000110_1_10_000_110_101_0_x_00;
      patterns[2285] = 32'b1011010100000110_1_11_000_110_101_0_x_00;
      patterns[2286] = 32'b0101010100000000_1_xx_000_xxx_101_0_1_01;
      patterns[2287] = 32'b0100010100000000_0_xx_000_101_xxx_1_x_xx;
      patterns[2288] = 32'b0000010110111101_1_xx_xxx_xxx_101_0_x_10;
      patterns[2289] = 32'b1000010100000111_1_00_000_111_101_0_x_00;
      patterns[2290] = 32'b1001010100000111_1_01_000_111_101_0_x_00;
      patterns[2291] = 32'b1010010100000111_1_10_000_111_101_0_x_00;
      patterns[2292] = 32'b1011010100000111_1_11_000_111_101_0_x_00;
      patterns[2293] = 32'b0101010100000000_1_xx_000_xxx_101_0_1_01;
      patterns[2294] = 32'b0100010100000000_0_xx_000_101_xxx_1_x_xx;
      patterns[2295] = 32'b0000010110001110_1_xx_xxx_xxx_101_0_x_10;
      patterns[2296] = 32'b1000010100010000_1_00_001_000_101_0_x_00;
      patterns[2297] = 32'b1001010100010000_1_01_001_000_101_0_x_00;
      patterns[2298] = 32'b1010010100010000_1_10_001_000_101_0_x_00;
      patterns[2299] = 32'b1011010100010000_1_11_001_000_101_0_x_00;
      patterns[2300] = 32'b0101010100010000_1_xx_001_xxx_101_0_1_01;
      patterns[2301] = 32'b0100010100010000_0_xx_001_101_xxx_1_x_xx;
      patterns[2302] = 32'b0000010100010100_1_xx_xxx_xxx_101_0_x_10;
      patterns[2303] = 32'b1000010100010001_1_00_001_001_101_0_x_00;
      patterns[2304] = 32'b1001010100010001_1_01_001_001_101_0_x_00;
      patterns[2305] = 32'b1010010100010001_1_10_001_001_101_0_x_00;
      patterns[2306] = 32'b1011010100010001_1_11_001_001_101_0_x_00;
      patterns[2307] = 32'b0101010100010000_1_xx_001_xxx_101_0_1_01;
      patterns[2308] = 32'b0100010100010000_0_xx_001_101_xxx_1_x_xx;
      patterns[2309] = 32'b0000010110101010_1_xx_xxx_xxx_101_0_x_10;
      patterns[2310] = 32'b1000010100010010_1_00_001_010_101_0_x_00;
      patterns[2311] = 32'b1001010100010010_1_01_001_010_101_0_x_00;
      patterns[2312] = 32'b1010010100010010_1_10_001_010_101_0_x_00;
      patterns[2313] = 32'b1011010100010010_1_11_001_010_101_0_x_00;
      patterns[2314] = 32'b0101010100010000_1_xx_001_xxx_101_0_1_01;
      patterns[2315] = 32'b0100010100010000_0_xx_001_101_xxx_1_x_xx;
      patterns[2316] = 32'b0000010101100110_1_xx_xxx_xxx_101_0_x_10;
      patterns[2317] = 32'b1000010100010011_1_00_001_011_101_0_x_00;
      patterns[2318] = 32'b1001010100010011_1_01_001_011_101_0_x_00;
      patterns[2319] = 32'b1010010100010011_1_10_001_011_101_0_x_00;
      patterns[2320] = 32'b1011010100010011_1_11_001_011_101_0_x_00;
      patterns[2321] = 32'b0101010100010000_1_xx_001_xxx_101_0_1_01;
      patterns[2322] = 32'b0100010100010000_0_xx_001_101_xxx_1_x_xx;
      patterns[2323] = 32'b0000010101011101_1_xx_xxx_xxx_101_0_x_10;
      patterns[2324] = 32'b1000010100010100_1_00_001_100_101_0_x_00;
      patterns[2325] = 32'b1001010100010100_1_01_001_100_101_0_x_00;
      patterns[2326] = 32'b1010010100010100_1_10_001_100_101_0_x_00;
      patterns[2327] = 32'b1011010100010100_1_11_001_100_101_0_x_00;
      patterns[2328] = 32'b0101010100010000_1_xx_001_xxx_101_0_1_01;
      patterns[2329] = 32'b0100010100010000_0_xx_001_101_xxx_1_x_xx;
      patterns[2330] = 32'b0000010100110000_1_xx_xxx_xxx_101_0_x_10;
      patterns[2331] = 32'b1000010100010101_1_00_001_101_101_0_x_00;
      patterns[2332] = 32'b1001010100010101_1_01_001_101_101_0_x_00;
      patterns[2333] = 32'b1010010100010101_1_10_001_101_101_0_x_00;
      patterns[2334] = 32'b1011010100010101_1_11_001_101_101_0_x_00;
      patterns[2335] = 32'b0101010100010000_1_xx_001_xxx_101_0_1_01;
      patterns[2336] = 32'b0100010100010000_0_xx_001_101_xxx_1_x_xx;
      patterns[2337] = 32'b0000010110001100_1_xx_xxx_xxx_101_0_x_10;
      patterns[2338] = 32'b1000010100010110_1_00_001_110_101_0_x_00;
      patterns[2339] = 32'b1001010100010110_1_01_001_110_101_0_x_00;
      patterns[2340] = 32'b1010010100010110_1_10_001_110_101_0_x_00;
      patterns[2341] = 32'b1011010100010110_1_11_001_110_101_0_x_00;
      patterns[2342] = 32'b0101010100010000_1_xx_001_xxx_101_0_1_01;
      patterns[2343] = 32'b0100010100010000_0_xx_001_101_xxx_1_x_xx;
      patterns[2344] = 32'b0000010101010101_1_xx_xxx_xxx_101_0_x_10;
      patterns[2345] = 32'b1000010100010111_1_00_001_111_101_0_x_00;
      patterns[2346] = 32'b1001010100010111_1_01_001_111_101_0_x_00;
      patterns[2347] = 32'b1010010100010111_1_10_001_111_101_0_x_00;
      patterns[2348] = 32'b1011010100010111_1_11_001_111_101_0_x_00;
      patterns[2349] = 32'b0101010100010000_1_xx_001_xxx_101_0_1_01;
      patterns[2350] = 32'b0100010100010000_0_xx_001_101_xxx_1_x_xx;
      patterns[2351] = 32'b0000010101001101_1_xx_xxx_xxx_101_0_x_10;
      patterns[2352] = 32'b1000010100100000_1_00_010_000_101_0_x_00;
      patterns[2353] = 32'b1001010100100000_1_01_010_000_101_0_x_00;
      patterns[2354] = 32'b1010010100100000_1_10_010_000_101_0_x_00;
      patterns[2355] = 32'b1011010100100000_1_11_010_000_101_0_x_00;
      patterns[2356] = 32'b0101010100100000_1_xx_010_xxx_101_0_1_01;
      patterns[2357] = 32'b0100010100100000_0_xx_010_101_xxx_1_x_xx;
      patterns[2358] = 32'b0000010100111000_1_xx_xxx_xxx_101_0_x_10;
      patterns[2359] = 32'b1000010100100001_1_00_010_001_101_0_x_00;
      patterns[2360] = 32'b1001010100100001_1_01_010_001_101_0_x_00;
      patterns[2361] = 32'b1010010100100001_1_10_010_001_101_0_x_00;
      patterns[2362] = 32'b1011010100100001_1_11_010_001_101_0_x_00;
      patterns[2363] = 32'b0101010100100000_1_xx_010_xxx_101_0_1_01;
      patterns[2364] = 32'b0100010100100000_0_xx_010_101_xxx_1_x_xx;
      patterns[2365] = 32'b0000010100001011_1_xx_xxx_xxx_101_0_x_10;
      patterns[2366] = 32'b1000010100100010_1_00_010_010_101_0_x_00;
      patterns[2367] = 32'b1001010100100010_1_01_010_010_101_0_x_00;
      patterns[2368] = 32'b1010010100100010_1_10_010_010_101_0_x_00;
      patterns[2369] = 32'b1011010100100010_1_11_010_010_101_0_x_00;
      patterns[2370] = 32'b0101010100100000_1_xx_010_xxx_101_0_1_01;
      patterns[2371] = 32'b0100010100100000_0_xx_010_101_xxx_1_x_xx;
      patterns[2372] = 32'b0000010101111011_1_xx_xxx_xxx_101_0_x_10;
      patterns[2373] = 32'b1000010100100011_1_00_010_011_101_0_x_00;
      patterns[2374] = 32'b1001010100100011_1_01_010_011_101_0_x_00;
      patterns[2375] = 32'b1010010100100011_1_10_010_011_101_0_x_00;
      patterns[2376] = 32'b1011010100100011_1_11_010_011_101_0_x_00;
      patterns[2377] = 32'b0101010100100000_1_xx_010_xxx_101_0_1_01;
      patterns[2378] = 32'b0100010100100000_0_xx_010_101_xxx_1_x_xx;
      patterns[2379] = 32'b0000010100011111_1_xx_xxx_xxx_101_0_x_10;
      patterns[2380] = 32'b1000010100100100_1_00_010_100_101_0_x_00;
      patterns[2381] = 32'b1001010100100100_1_01_010_100_101_0_x_00;
      patterns[2382] = 32'b1010010100100100_1_10_010_100_101_0_x_00;
      patterns[2383] = 32'b1011010100100100_1_11_010_100_101_0_x_00;
      patterns[2384] = 32'b0101010100100000_1_xx_010_xxx_101_0_1_01;
      patterns[2385] = 32'b0100010100100000_0_xx_010_101_xxx_1_x_xx;
      patterns[2386] = 32'b0000010101111110_1_xx_xxx_xxx_101_0_x_10;
      patterns[2387] = 32'b1000010100100101_1_00_010_101_101_0_x_00;
      patterns[2388] = 32'b1001010100100101_1_01_010_101_101_0_x_00;
      patterns[2389] = 32'b1010010100100101_1_10_010_101_101_0_x_00;
      patterns[2390] = 32'b1011010100100101_1_11_010_101_101_0_x_00;
      patterns[2391] = 32'b0101010100100000_1_xx_010_xxx_101_0_1_01;
      patterns[2392] = 32'b0100010100100000_0_xx_010_101_xxx_1_x_xx;
      patterns[2393] = 32'b0000010100001111_1_xx_xxx_xxx_101_0_x_10;
      patterns[2394] = 32'b1000010100100110_1_00_010_110_101_0_x_00;
      patterns[2395] = 32'b1001010100100110_1_01_010_110_101_0_x_00;
      patterns[2396] = 32'b1010010100100110_1_10_010_110_101_0_x_00;
      patterns[2397] = 32'b1011010100100110_1_11_010_110_101_0_x_00;
      patterns[2398] = 32'b0101010100100000_1_xx_010_xxx_101_0_1_01;
      patterns[2399] = 32'b0100010100100000_0_xx_010_101_xxx_1_x_xx;
      patterns[2400] = 32'b0000010111100001_1_xx_xxx_xxx_101_0_x_10;
      patterns[2401] = 32'b1000010100100111_1_00_010_111_101_0_x_00;
      patterns[2402] = 32'b1001010100100111_1_01_010_111_101_0_x_00;
      patterns[2403] = 32'b1010010100100111_1_10_010_111_101_0_x_00;
      patterns[2404] = 32'b1011010100100111_1_11_010_111_101_0_x_00;
      patterns[2405] = 32'b0101010100100000_1_xx_010_xxx_101_0_1_01;
      patterns[2406] = 32'b0100010100100000_0_xx_010_101_xxx_1_x_xx;
      patterns[2407] = 32'b0000010110000001_1_xx_xxx_xxx_101_0_x_10;
      patterns[2408] = 32'b1000010100110000_1_00_011_000_101_0_x_00;
      patterns[2409] = 32'b1001010100110000_1_01_011_000_101_0_x_00;
      patterns[2410] = 32'b1010010100110000_1_10_011_000_101_0_x_00;
      patterns[2411] = 32'b1011010100110000_1_11_011_000_101_0_x_00;
      patterns[2412] = 32'b0101010100110000_1_xx_011_xxx_101_0_1_01;
      patterns[2413] = 32'b0100010100110000_0_xx_011_101_xxx_1_x_xx;
      patterns[2414] = 32'b0000010111001111_1_xx_xxx_xxx_101_0_x_10;
      patterns[2415] = 32'b1000010100110001_1_00_011_001_101_0_x_00;
      patterns[2416] = 32'b1001010100110001_1_01_011_001_101_0_x_00;
      patterns[2417] = 32'b1010010100110001_1_10_011_001_101_0_x_00;
      patterns[2418] = 32'b1011010100110001_1_11_011_001_101_0_x_00;
      patterns[2419] = 32'b0101010100110000_1_xx_011_xxx_101_0_1_01;
      patterns[2420] = 32'b0100010100110000_0_xx_011_101_xxx_1_x_xx;
      patterns[2421] = 32'b0000010101110001_1_xx_xxx_xxx_101_0_x_10;
      patterns[2422] = 32'b1000010100110010_1_00_011_010_101_0_x_00;
      patterns[2423] = 32'b1001010100110010_1_01_011_010_101_0_x_00;
      patterns[2424] = 32'b1010010100110010_1_10_011_010_101_0_x_00;
      patterns[2425] = 32'b1011010100110010_1_11_011_010_101_0_x_00;
      patterns[2426] = 32'b0101010100110000_1_xx_011_xxx_101_0_1_01;
      patterns[2427] = 32'b0100010100110000_0_xx_011_101_xxx_1_x_xx;
      patterns[2428] = 32'b0000010110110111_1_xx_xxx_xxx_101_0_x_10;
      patterns[2429] = 32'b1000010100110011_1_00_011_011_101_0_x_00;
      patterns[2430] = 32'b1001010100110011_1_01_011_011_101_0_x_00;
      patterns[2431] = 32'b1010010100110011_1_10_011_011_101_0_x_00;
      patterns[2432] = 32'b1011010100110011_1_11_011_011_101_0_x_00;
      patterns[2433] = 32'b0101010100110000_1_xx_011_xxx_101_0_1_01;
      patterns[2434] = 32'b0100010100110000_0_xx_011_101_xxx_1_x_xx;
      patterns[2435] = 32'b0000010110100110_1_xx_xxx_xxx_101_0_x_10;
      patterns[2436] = 32'b1000010100110100_1_00_011_100_101_0_x_00;
      patterns[2437] = 32'b1001010100110100_1_01_011_100_101_0_x_00;
      patterns[2438] = 32'b1010010100110100_1_10_011_100_101_0_x_00;
      patterns[2439] = 32'b1011010100110100_1_11_011_100_101_0_x_00;
      patterns[2440] = 32'b0101010100110000_1_xx_011_xxx_101_0_1_01;
      patterns[2441] = 32'b0100010100110000_0_xx_011_101_xxx_1_x_xx;
      patterns[2442] = 32'b0000010100111110_1_xx_xxx_xxx_101_0_x_10;
      patterns[2443] = 32'b1000010100110101_1_00_011_101_101_0_x_00;
      patterns[2444] = 32'b1001010100110101_1_01_011_101_101_0_x_00;
      patterns[2445] = 32'b1010010100110101_1_10_011_101_101_0_x_00;
      patterns[2446] = 32'b1011010100110101_1_11_011_101_101_0_x_00;
      patterns[2447] = 32'b0101010100110000_1_xx_011_xxx_101_0_1_01;
      patterns[2448] = 32'b0100010100110000_0_xx_011_101_xxx_1_x_xx;
      patterns[2449] = 32'b0000010111111010_1_xx_xxx_xxx_101_0_x_10;
      patterns[2450] = 32'b1000010100110110_1_00_011_110_101_0_x_00;
      patterns[2451] = 32'b1001010100110110_1_01_011_110_101_0_x_00;
      patterns[2452] = 32'b1010010100110110_1_10_011_110_101_0_x_00;
      patterns[2453] = 32'b1011010100110110_1_11_011_110_101_0_x_00;
      patterns[2454] = 32'b0101010100110000_1_xx_011_xxx_101_0_1_01;
      patterns[2455] = 32'b0100010100110000_0_xx_011_101_xxx_1_x_xx;
      patterns[2456] = 32'b0000010111011000_1_xx_xxx_xxx_101_0_x_10;
      patterns[2457] = 32'b1000010100110111_1_00_011_111_101_0_x_00;
      patterns[2458] = 32'b1001010100110111_1_01_011_111_101_0_x_00;
      patterns[2459] = 32'b1010010100110111_1_10_011_111_101_0_x_00;
      patterns[2460] = 32'b1011010100110111_1_11_011_111_101_0_x_00;
      patterns[2461] = 32'b0101010100110000_1_xx_011_xxx_101_0_1_01;
      patterns[2462] = 32'b0100010100110000_0_xx_011_101_xxx_1_x_xx;
      patterns[2463] = 32'b0000010100001111_1_xx_xxx_xxx_101_0_x_10;
      patterns[2464] = 32'b1000010101000000_1_00_100_000_101_0_x_00;
      patterns[2465] = 32'b1001010101000000_1_01_100_000_101_0_x_00;
      patterns[2466] = 32'b1010010101000000_1_10_100_000_101_0_x_00;
      patterns[2467] = 32'b1011010101000000_1_11_100_000_101_0_x_00;
      patterns[2468] = 32'b0101010101000000_1_xx_100_xxx_101_0_1_01;
      patterns[2469] = 32'b0100010101000000_0_xx_100_101_xxx_1_x_xx;
      patterns[2470] = 32'b0000010111100110_1_xx_xxx_xxx_101_0_x_10;
      patterns[2471] = 32'b1000010101000001_1_00_100_001_101_0_x_00;
      patterns[2472] = 32'b1001010101000001_1_01_100_001_101_0_x_00;
      patterns[2473] = 32'b1010010101000001_1_10_100_001_101_0_x_00;
      patterns[2474] = 32'b1011010101000001_1_11_100_001_101_0_x_00;
      patterns[2475] = 32'b0101010101000000_1_xx_100_xxx_101_0_1_01;
      patterns[2476] = 32'b0100010101000000_0_xx_100_101_xxx_1_x_xx;
      patterns[2477] = 32'b0000010100110001_1_xx_xxx_xxx_101_0_x_10;
      patterns[2478] = 32'b1000010101000010_1_00_100_010_101_0_x_00;
      patterns[2479] = 32'b1001010101000010_1_01_100_010_101_0_x_00;
      patterns[2480] = 32'b1010010101000010_1_10_100_010_101_0_x_00;
      patterns[2481] = 32'b1011010101000010_1_11_100_010_101_0_x_00;
      patterns[2482] = 32'b0101010101000000_1_xx_100_xxx_101_0_1_01;
      patterns[2483] = 32'b0100010101000000_0_xx_100_101_xxx_1_x_xx;
      patterns[2484] = 32'b0000010111000110_1_xx_xxx_xxx_101_0_x_10;
      patterns[2485] = 32'b1000010101000011_1_00_100_011_101_0_x_00;
      patterns[2486] = 32'b1001010101000011_1_01_100_011_101_0_x_00;
      patterns[2487] = 32'b1010010101000011_1_10_100_011_101_0_x_00;
      patterns[2488] = 32'b1011010101000011_1_11_100_011_101_0_x_00;
      patterns[2489] = 32'b0101010101000000_1_xx_100_xxx_101_0_1_01;
      patterns[2490] = 32'b0100010101000000_0_xx_100_101_xxx_1_x_xx;
      patterns[2491] = 32'b0000010101110100_1_xx_xxx_xxx_101_0_x_10;
      patterns[2492] = 32'b1000010101000100_1_00_100_100_101_0_x_00;
      patterns[2493] = 32'b1001010101000100_1_01_100_100_101_0_x_00;
      patterns[2494] = 32'b1010010101000100_1_10_100_100_101_0_x_00;
      patterns[2495] = 32'b1011010101000100_1_11_100_100_101_0_x_00;
      patterns[2496] = 32'b0101010101000000_1_xx_100_xxx_101_0_1_01;
      patterns[2497] = 32'b0100010101000000_0_xx_100_101_xxx_1_x_xx;
      patterns[2498] = 32'b0000010110000000_1_xx_xxx_xxx_101_0_x_10;
      patterns[2499] = 32'b1000010101000101_1_00_100_101_101_0_x_00;
      patterns[2500] = 32'b1001010101000101_1_01_100_101_101_0_x_00;
      patterns[2501] = 32'b1010010101000101_1_10_100_101_101_0_x_00;
      patterns[2502] = 32'b1011010101000101_1_11_100_101_101_0_x_00;
      patterns[2503] = 32'b0101010101000000_1_xx_100_xxx_101_0_1_01;
      patterns[2504] = 32'b0100010101000000_0_xx_100_101_xxx_1_x_xx;
      patterns[2505] = 32'b0000010111010000_1_xx_xxx_xxx_101_0_x_10;
      patterns[2506] = 32'b1000010101000110_1_00_100_110_101_0_x_00;
      patterns[2507] = 32'b1001010101000110_1_01_100_110_101_0_x_00;
      patterns[2508] = 32'b1010010101000110_1_10_100_110_101_0_x_00;
      patterns[2509] = 32'b1011010101000110_1_11_100_110_101_0_x_00;
      patterns[2510] = 32'b0101010101000000_1_xx_100_xxx_101_0_1_01;
      patterns[2511] = 32'b0100010101000000_0_xx_100_101_xxx_1_x_xx;
      patterns[2512] = 32'b0000010100101000_1_xx_xxx_xxx_101_0_x_10;
      patterns[2513] = 32'b1000010101000111_1_00_100_111_101_0_x_00;
      patterns[2514] = 32'b1001010101000111_1_01_100_111_101_0_x_00;
      patterns[2515] = 32'b1010010101000111_1_10_100_111_101_0_x_00;
      patterns[2516] = 32'b1011010101000111_1_11_100_111_101_0_x_00;
      patterns[2517] = 32'b0101010101000000_1_xx_100_xxx_101_0_1_01;
      patterns[2518] = 32'b0100010101000000_0_xx_100_101_xxx_1_x_xx;
      patterns[2519] = 32'b0000010111110101_1_xx_xxx_xxx_101_0_x_10;
      patterns[2520] = 32'b1000010101010000_1_00_101_000_101_0_x_00;
      patterns[2521] = 32'b1001010101010000_1_01_101_000_101_0_x_00;
      patterns[2522] = 32'b1010010101010000_1_10_101_000_101_0_x_00;
      patterns[2523] = 32'b1011010101010000_1_11_101_000_101_0_x_00;
      patterns[2524] = 32'b0101010101010000_1_xx_101_xxx_101_0_1_01;
      patterns[2525] = 32'b0100010101010000_0_xx_101_101_xxx_1_x_xx;
      patterns[2526] = 32'b0000010111011011_1_xx_xxx_xxx_101_0_x_10;
      patterns[2527] = 32'b1000010101010001_1_00_101_001_101_0_x_00;
      patterns[2528] = 32'b1001010101010001_1_01_101_001_101_0_x_00;
      patterns[2529] = 32'b1010010101010001_1_10_101_001_101_0_x_00;
      patterns[2530] = 32'b1011010101010001_1_11_101_001_101_0_x_00;
      patterns[2531] = 32'b0101010101010000_1_xx_101_xxx_101_0_1_01;
      patterns[2532] = 32'b0100010101010000_0_xx_101_101_xxx_1_x_xx;
      patterns[2533] = 32'b0000010101101000_1_xx_xxx_xxx_101_0_x_10;
      patterns[2534] = 32'b1000010101010010_1_00_101_010_101_0_x_00;
      patterns[2535] = 32'b1001010101010010_1_01_101_010_101_0_x_00;
      patterns[2536] = 32'b1010010101010010_1_10_101_010_101_0_x_00;
      patterns[2537] = 32'b1011010101010010_1_11_101_010_101_0_x_00;
      patterns[2538] = 32'b0101010101010000_1_xx_101_xxx_101_0_1_01;
      patterns[2539] = 32'b0100010101010000_0_xx_101_101_xxx_1_x_xx;
      patterns[2540] = 32'b0000010101101000_1_xx_xxx_xxx_101_0_x_10;
      patterns[2541] = 32'b1000010101010011_1_00_101_011_101_0_x_00;
      patterns[2542] = 32'b1001010101010011_1_01_101_011_101_0_x_00;
      patterns[2543] = 32'b1010010101010011_1_10_101_011_101_0_x_00;
      patterns[2544] = 32'b1011010101010011_1_11_101_011_101_0_x_00;
      patterns[2545] = 32'b0101010101010000_1_xx_101_xxx_101_0_1_01;
      patterns[2546] = 32'b0100010101010000_0_xx_101_101_xxx_1_x_xx;
      patterns[2547] = 32'b0000010100010111_1_xx_xxx_xxx_101_0_x_10;
      patterns[2548] = 32'b1000010101010100_1_00_101_100_101_0_x_00;
      patterns[2549] = 32'b1001010101010100_1_01_101_100_101_0_x_00;
      patterns[2550] = 32'b1010010101010100_1_10_101_100_101_0_x_00;
      patterns[2551] = 32'b1011010101010100_1_11_101_100_101_0_x_00;
      patterns[2552] = 32'b0101010101010000_1_xx_101_xxx_101_0_1_01;
      patterns[2553] = 32'b0100010101010000_0_xx_101_101_xxx_1_x_xx;
      patterns[2554] = 32'b0000010101110100_1_xx_xxx_xxx_101_0_x_10;
      patterns[2555] = 32'b1000010101010101_1_00_101_101_101_0_x_00;
      patterns[2556] = 32'b1001010101010101_1_01_101_101_101_0_x_00;
      patterns[2557] = 32'b1010010101010101_1_10_101_101_101_0_x_00;
      patterns[2558] = 32'b1011010101010101_1_11_101_101_101_0_x_00;
      patterns[2559] = 32'b0101010101010000_1_xx_101_xxx_101_0_1_01;
      patterns[2560] = 32'b0100010101010000_0_xx_101_101_xxx_1_x_xx;
      patterns[2561] = 32'b0000010111011011_1_xx_xxx_xxx_101_0_x_10;
      patterns[2562] = 32'b1000010101010110_1_00_101_110_101_0_x_00;
      patterns[2563] = 32'b1001010101010110_1_01_101_110_101_0_x_00;
      patterns[2564] = 32'b1010010101010110_1_10_101_110_101_0_x_00;
      patterns[2565] = 32'b1011010101010110_1_11_101_110_101_0_x_00;
      patterns[2566] = 32'b0101010101010000_1_xx_101_xxx_101_0_1_01;
      patterns[2567] = 32'b0100010101010000_0_xx_101_101_xxx_1_x_xx;
      patterns[2568] = 32'b0000010100011011_1_xx_xxx_xxx_101_0_x_10;
      patterns[2569] = 32'b1000010101010111_1_00_101_111_101_0_x_00;
      patterns[2570] = 32'b1001010101010111_1_01_101_111_101_0_x_00;
      patterns[2571] = 32'b1010010101010111_1_10_101_111_101_0_x_00;
      patterns[2572] = 32'b1011010101010111_1_11_101_111_101_0_x_00;
      patterns[2573] = 32'b0101010101010000_1_xx_101_xxx_101_0_1_01;
      patterns[2574] = 32'b0100010101010000_0_xx_101_101_xxx_1_x_xx;
      patterns[2575] = 32'b0000010100100111_1_xx_xxx_xxx_101_0_x_10;
      patterns[2576] = 32'b1000010101100000_1_00_110_000_101_0_x_00;
      patterns[2577] = 32'b1001010101100000_1_01_110_000_101_0_x_00;
      patterns[2578] = 32'b1010010101100000_1_10_110_000_101_0_x_00;
      patterns[2579] = 32'b1011010101100000_1_11_110_000_101_0_x_00;
      patterns[2580] = 32'b0101010101100000_1_xx_110_xxx_101_0_1_01;
      patterns[2581] = 32'b0100010101100000_0_xx_110_101_xxx_1_x_xx;
      patterns[2582] = 32'b0000010111100010_1_xx_xxx_xxx_101_0_x_10;
      patterns[2583] = 32'b1000010101100001_1_00_110_001_101_0_x_00;
      patterns[2584] = 32'b1001010101100001_1_01_110_001_101_0_x_00;
      patterns[2585] = 32'b1010010101100001_1_10_110_001_101_0_x_00;
      patterns[2586] = 32'b1011010101100001_1_11_110_001_101_0_x_00;
      patterns[2587] = 32'b0101010101100000_1_xx_110_xxx_101_0_1_01;
      patterns[2588] = 32'b0100010101100000_0_xx_110_101_xxx_1_x_xx;
      patterns[2589] = 32'b0000010111000110_1_xx_xxx_xxx_101_0_x_10;
      patterns[2590] = 32'b1000010101100010_1_00_110_010_101_0_x_00;
      patterns[2591] = 32'b1001010101100010_1_01_110_010_101_0_x_00;
      patterns[2592] = 32'b1010010101100010_1_10_110_010_101_0_x_00;
      patterns[2593] = 32'b1011010101100010_1_11_110_010_101_0_x_00;
      patterns[2594] = 32'b0101010101100000_1_xx_110_xxx_101_0_1_01;
      patterns[2595] = 32'b0100010101100000_0_xx_110_101_xxx_1_x_xx;
      patterns[2596] = 32'b0000010111110110_1_xx_xxx_xxx_101_0_x_10;
      patterns[2597] = 32'b1000010101100011_1_00_110_011_101_0_x_00;
      patterns[2598] = 32'b1001010101100011_1_01_110_011_101_0_x_00;
      patterns[2599] = 32'b1010010101100011_1_10_110_011_101_0_x_00;
      patterns[2600] = 32'b1011010101100011_1_11_110_011_101_0_x_00;
      patterns[2601] = 32'b0101010101100000_1_xx_110_xxx_101_0_1_01;
      patterns[2602] = 32'b0100010101100000_0_xx_110_101_xxx_1_x_xx;
      patterns[2603] = 32'b0000010110111011_1_xx_xxx_xxx_101_0_x_10;
      patterns[2604] = 32'b1000010101100100_1_00_110_100_101_0_x_00;
      patterns[2605] = 32'b1001010101100100_1_01_110_100_101_0_x_00;
      patterns[2606] = 32'b1010010101100100_1_10_110_100_101_0_x_00;
      patterns[2607] = 32'b1011010101100100_1_11_110_100_101_0_x_00;
      patterns[2608] = 32'b0101010101100000_1_xx_110_xxx_101_0_1_01;
      patterns[2609] = 32'b0100010101100000_0_xx_110_101_xxx_1_x_xx;
      patterns[2610] = 32'b0000010101100001_1_xx_xxx_xxx_101_0_x_10;
      patterns[2611] = 32'b1000010101100101_1_00_110_101_101_0_x_00;
      patterns[2612] = 32'b1001010101100101_1_01_110_101_101_0_x_00;
      patterns[2613] = 32'b1010010101100101_1_10_110_101_101_0_x_00;
      patterns[2614] = 32'b1011010101100101_1_11_110_101_101_0_x_00;
      patterns[2615] = 32'b0101010101100000_1_xx_110_xxx_101_0_1_01;
      patterns[2616] = 32'b0100010101100000_0_xx_110_101_xxx_1_x_xx;
      patterns[2617] = 32'b0000010111010110_1_xx_xxx_xxx_101_0_x_10;
      patterns[2618] = 32'b1000010101100110_1_00_110_110_101_0_x_00;
      patterns[2619] = 32'b1001010101100110_1_01_110_110_101_0_x_00;
      patterns[2620] = 32'b1010010101100110_1_10_110_110_101_0_x_00;
      patterns[2621] = 32'b1011010101100110_1_11_110_110_101_0_x_00;
      patterns[2622] = 32'b0101010101100000_1_xx_110_xxx_101_0_1_01;
      patterns[2623] = 32'b0100010101100000_0_xx_110_101_xxx_1_x_xx;
      patterns[2624] = 32'b0000010101101101_1_xx_xxx_xxx_101_0_x_10;
      patterns[2625] = 32'b1000010101100111_1_00_110_111_101_0_x_00;
      patterns[2626] = 32'b1001010101100111_1_01_110_111_101_0_x_00;
      patterns[2627] = 32'b1010010101100111_1_10_110_111_101_0_x_00;
      patterns[2628] = 32'b1011010101100111_1_11_110_111_101_0_x_00;
      patterns[2629] = 32'b0101010101100000_1_xx_110_xxx_101_0_1_01;
      patterns[2630] = 32'b0100010101100000_0_xx_110_101_xxx_1_x_xx;
      patterns[2631] = 32'b0000010111110011_1_xx_xxx_xxx_101_0_x_10;
      patterns[2632] = 32'b1000010101110000_1_00_111_000_101_0_x_00;
      patterns[2633] = 32'b1001010101110000_1_01_111_000_101_0_x_00;
      patterns[2634] = 32'b1010010101110000_1_10_111_000_101_0_x_00;
      patterns[2635] = 32'b1011010101110000_1_11_111_000_101_0_x_00;
      patterns[2636] = 32'b0101010101110000_1_xx_111_xxx_101_0_1_01;
      patterns[2637] = 32'b0100010101110000_0_xx_111_101_xxx_1_x_xx;
      patterns[2638] = 32'b0000010101110011_1_xx_xxx_xxx_101_0_x_10;
      patterns[2639] = 32'b1000010101110001_1_00_111_001_101_0_x_00;
      patterns[2640] = 32'b1001010101110001_1_01_111_001_101_0_x_00;
      patterns[2641] = 32'b1010010101110001_1_10_111_001_101_0_x_00;
      patterns[2642] = 32'b1011010101110001_1_11_111_001_101_0_x_00;
      patterns[2643] = 32'b0101010101110000_1_xx_111_xxx_101_0_1_01;
      patterns[2644] = 32'b0100010101110000_0_xx_111_101_xxx_1_x_xx;
      patterns[2645] = 32'b0000010101100101_1_xx_xxx_xxx_101_0_x_10;
      patterns[2646] = 32'b1000010101110010_1_00_111_010_101_0_x_00;
      patterns[2647] = 32'b1001010101110010_1_01_111_010_101_0_x_00;
      patterns[2648] = 32'b1010010101110010_1_10_111_010_101_0_x_00;
      patterns[2649] = 32'b1011010101110010_1_11_111_010_101_0_x_00;
      patterns[2650] = 32'b0101010101110000_1_xx_111_xxx_101_0_1_01;
      patterns[2651] = 32'b0100010101110000_0_xx_111_101_xxx_1_x_xx;
      patterns[2652] = 32'b0000010101011110_1_xx_xxx_xxx_101_0_x_10;
      patterns[2653] = 32'b1000010101110011_1_00_111_011_101_0_x_00;
      patterns[2654] = 32'b1001010101110011_1_01_111_011_101_0_x_00;
      patterns[2655] = 32'b1010010101110011_1_10_111_011_101_0_x_00;
      patterns[2656] = 32'b1011010101110011_1_11_111_011_101_0_x_00;
      patterns[2657] = 32'b0101010101110000_1_xx_111_xxx_101_0_1_01;
      patterns[2658] = 32'b0100010101110000_0_xx_111_101_xxx_1_x_xx;
      patterns[2659] = 32'b0000010100011001_1_xx_xxx_xxx_101_0_x_10;
      patterns[2660] = 32'b1000010101110100_1_00_111_100_101_0_x_00;
      patterns[2661] = 32'b1001010101110100_1_01_111_100_101_0_x_00;
      patterns[2662] = 32'b1010010101110100_1_10_111_100_101_0_x_00;
      patterns[2663] = 32'b1011010101110100_1_11_111_100_101_0_x_00;
      patterns[2664] = 32'b0101010101110000_1_xx_111_xxx_101_0_1_01;
      patterns[2665] = 32'b0100010101110000_0_xx_111_101_xxx_1_x_xx;
      patterns[2666] = 32'b0000010110000101_1_xx_xxx_xxx_101_0_x_10;
      patterns[2667] = 32'b1000010101110101_1_00_111_101_101_0_x_00;
      patterns[2668] = 32'b1001010101110101_1_01_111_101_101_0_x_00;
      patterns[2669] = 32'b1010010101110101_1_10_111_101_101_0_x_00;
      patterns[2670] = 32'b1011010101110101_1_11_111_101_101_0_x_00;
      patterns[2671] = 32'b0101010101110000_1_xx_111_xxx_101_0_1_01;
      patterns[2672] = 32'b0100010101110000_0_xx_111_101_xxx_1_x_xx;
      patterns[2673] = 32'b0000010101011001_1_xx_xxx_xxx_101_0_x_10;
      patterns[2674] = 32'b1000010101110110_1_00_111_110_101_0_x_00;
      patterns[2675] = 32'b1001010101110110_1_01_111_110_101_0_x_00;
      patterns[2676] = 32'b1010010101110110_1_10_111_110_101_0_x_00;
      patterns[2677] = 32'b1011010101110110_1_11_111_110_101_0_x_00;
      patterns[2678] = 32'b0101010101110000_1_xx_111_xxx_101_0_1_01;
      patterns[2679] = 32'b0100010101110000_0_xx_111_101_xxx_1_x_xx;
      patterns[2680] = 32'b0000010111111100_1_xx_xxx_xxx_101_0_x_10;
      patterns[2681] = 32'b1000010101110111_1_00_111_111_101_0_x_00;
      patterns[2682] = 32'b1001010101110111_1_01_111_111_101_0_x_00;
      patterns[2683] = 32'b1010010101110111_1_10_111_111_101_0_x_00;
      patterns[2684] = 32'b1011010101110111_1_11_111_111_101_0_x_00;
      patterns[2685] = 32'b0101010101110000_1_xx_111_xxx_101_0_1_01;
      patterns[2686] = 32'b0100010101110000_0_xx_111_101_xxx_1_x_xx;
      patterns[2687] = 32'b0000010111100000_1_xx_xxx_xxx_101_0_x_10;
      patterns[2688] = 32'b1000011000000000_1_00_000_000_110_0_x_00;
      patterns[2689] = 32'b1001011000000000_1_01_000_000_110_0_x_00;
      patterns[2690] = 32'b1010011000000000_1_10_000_000_110_0_x_00;
      patterns[2691] = 32'b1011011000000000_1_11_000_000_110_0_x_00;
      patterns[2692] = 32'b0101011000000000_1_xx_000_xxx_110_0_1_01;
      patterns[2693] = 32'b0100011000000000_0_xx_000_110_xxx_1_x_xx;
      patterns[2694] = 32'b0000011001111110_1_xx_xxx_xxx_110_0_x_10;
      patterns[2695] = 32'b1000011000000001_1_00_000_001_110_0_x_00;
      patterns[2696] = 32'b1001011000000001_1_01_000_001_110_0_x_00;
      patterns[2697] = 32'b1010011000000001_1_10_000_001_110_0_x_00;
      patterns[2698] = 32'b1011011000000001_1_11_000_001_110_0_x_00;
      patterns[2699] = 32'b0101011000000000_1_xx_000_xxx_110_0_1_01;
      patterns[2700] = 32'b0100011000000000_0_xx_000_110_xxx_1_x_xx;
      patterns[2701] = 32'b0000011001101100_1_xx_xxx_xxx_110_0_x_10;
      patterns[2702] = 32'b1000011000000010_1_00_000_010_110_0_x_00;
      patterns[2703] = 32'b1001011000000010_1_01_000_010_110_0_x_00;
      patterns[2704] = 32'b1010011000000010_1_10_000_010_110_0_x_00;
      patterns[2705] = 32'b1011011000000010_1_11_000_010_110_0_x_00;
      patterns[2706] = 32'b0101011000000000_1_xx_000_xxx_110_0_1_01;
      patterns[2707] = 32'b0100011000000000_0_xx_000_110_xxx_1_x_xx;
      patterns[2708] = 32'b0000011010101111_1_xx_xxx_xxx_110_0_x_10;
      patterns[2709] = 32'b1000011000000011_1_00_000_011_110_0_x_00;
      patterns[2710] = 32'b1001011000000011_1_01_000_011_110_0_x_00;
      patterns[2711] = 32'b1010011000000011_1_10_000_011_110_0_x_00;
      patterns[2712] = 32'b1011011000000011_1_11_000_011_110_0_x_00;
      patterns[2713] = 32'b0101011000000000_1_xx_000_xxx_110_0_1_01;
      patterns[2714] = 32'b0100011000000000_0_xx_000_110_xxx_1_x_xx;
      patterns[2715] = 32'b0000011001011110_1_xx_xxx_xxx_110_0_x_10;
      patterns[2716] = 32'b1000011000000100_1_00_000_100_110_0_x_00;
      patterns[2717] = 32'b1001011000000100_1_01_000_100_110_0_x_00;
      patterns[2718] = 32'b1010011000000100_1_10_000_100_110_0_x_00;
      patterns[2719] = 32'b1011011000000100_1_11_000_100_110_0_x_00;
      patterns[2720] = 32'b0101011000000000_1_xx_000_xxx_110_0_1_01;
      patterns[2721] = 32'b0100011000000000_0_xx_000_110_xxx_1_x_xx;
      patterns[2722] = 32'b0000011001011001_1_xx_xxx_xxx_110_0_x_10;
      patterns[2723] = 32'b1000011000000101_1_00_000_101_110_0_x_00;
      patterns[2724] = 32'b1001011000000101_1_01_000_101_110_0_x_00;
      patterns[2725] = 32'b1010011000000101_1_10_000_101_110_0_x_00;
      patterns[2726] = 32'b1011011000000101_1_11_000_101_110_0_x_00;
      patterns[2727] = 32'b0101011000000000_1_xx_000_xxx_110_0_1_01;
      patterns[2728] = 32'b0100011000000000_0_xx_000_110_xxx_1_x_xx;
      patterns[2729] = 32'b0000011010000000_1_xx_xxx_xxx_110_0_x_10;
      patterns[2730] = 32'b1000011000000110_1_00_000_110_110_0_x_00;
      patterns[2731] = 32'b1001011000000110_1_01_000_110_110_0_x_00;
      patterns[2732] = 32'b1010011000000110_1_10_000_110_110_0_x_00;
      patterns[2733] = 32'b1011011000000110_1_11_000_110_110_0_x_00;
      patterns[2734] = 32'b0101011000000000_1_xx_000_xxx_110_0_1_01;
      patterns[2735] = 32'b0100011000000000_0_xx_000_110_xxx_1_x_xx;
      patterns[2736] = 32'b0000011011000101_1_xx_xxx_xxx_110_0_x_10;
      patterns[2737] = 32'b1000011000000111_1_00_000_111_110_0_x_00;
      patterns[2738] = 32'b1001011000000111_1_01_000_111_110_0_x_00;
      patterns[2739] = 32'b1010011000000111_1_10_000_111_110_0_x_00;
      patterns[2740] = 32'b1011011000000111_1_11_000_111_110_0_x_00;
      patterns[2741] = 32'b0101011000000000_1_xx_000_xxx_110_0_1_01;
      patterns[2742] = 32'b0100011000000000_0_xx_000_110_xxx_1_x_xx;
      patterns[2743] = 32'b0000011001010011_1_xx_xxx_xxx_110_0_x_10;
      patterns[2744] = 32'b1000011000010000_1_00_001_000_110_0_x_00;
      patterns[2745] = 32'b1001011000010000_1_01_001_000_110_0_x_00;
      patterns[2746] = 32'b1010011000010000_1_10_001_000_110_0_x_00;
      patterns[2747] = 32'b1011011000010000_1_11_001_000_110_0_x_00;
      patterns[2748] = 32'b0101011000010000_1_xx_001_xxx_110_0_1_01;
      patterns[2749] = 32'b0100011000010000_0_xx_001_110_xxx_1_x_xx;
      patterns[2750] = 32'b0000011001011011_1_xx_xxx_xxx_110_0_x_10;
      patterns[2751] = 32'b1000011000010001_1_00_001_001_110_0_x_00;
      patterns[2752] = 32'b1001011000010001_1_01_001_001_110_0_x_00;
      patterns[2753] = 32'b1010011000010001_1_10_001_001_110_0_x_00;
      patterns[2754] = 32'b1011011000010001_1_11_001_001_110_0_x_00;
      patterns[2755] = 32'b0101011000010000_1_xx_001_xxx_110_0_1_01;
      patterns[2756] = 32'b0100011000010000_0_xx_001_110_xxx_1_x_xx;
      patterns[2757] = 32'b0000011010011011_1_xx_xxx_xxx_110_0_x_10;
      patterns[2758] = 32'b1000011000010010_1_00_001_010_110_0_x_00;
      patterns[2759] = 32'b1001011000010010_1_01_001_010_110_0_x_00;
      patterns[2760] = 32'b1010011000010010_1_10_001_010_110_0_x_00;
      patterns[2761] = 32'b1011011000010010_1_11_001_010_110_0_x_00;
      patterns[2762] = 32'b0101011000010000_1_xx_001_xxx_110_0_1_01;
      patterns[2763] = 32'b0100011000010000_0_xx_001_110_xxx_1_x_xx;
      patterns[2764] = 32'b0000011010010010_1_xx_xxx_xxx_110_0_x_10;
      patterns[2765] = 32'b1000011000010011_1_00_001_011_110_0_x_00;
      patterns[2766] = 32'b1001011000010011_1_01_001_011_110_0_x_00;
      patterns[2767] = 32'b1010011000010011_1_10_001_011_110_0_x_00;
      patterns[2768] = 32'b1011011000010011_1_11_001_011_110_0_x_00;
      patterns[2769] = 32'b0101011000010000_1_xx_001_xxx_110_0_1_01;
      patterns[2770] = 32'b0100011000010000_0_xx_001_110_xxx_1_x_xx;
      patterns[2771] = 32'b0000011011101001_1_xx_xxx_xxx_110_0_x_10;
      patterns[2772] = 32'b1000011000010100_1_00_001_100_110_0_x_00;
      patterns[2773] = 32'b1001011000010100_1_01_001_100_110_0_x_00;
      patterns[2774] = 32'b1010011000010100_1_10_001_100_110_0_x_00;
      patterns[2775] = 32'b1011011000010100_1_11_001_100_110_0_x_00;
      patterns[2776] = 32'b0101011000010000_1_xx_001_xxx_110_0_1_01;
      patterns[2777] = 32'b0100011000010000_0_xx_001_110_xxx_1_x_xx;
      patterns[2778] = 32'b0000011011000011_1_xx_xxx_xxx_110_0_x_10;
      patterns[2779] = 32'b1000011000010101_1_00_001_101_110_0_x_00;
      patterns[2780] = 32'b1001011000010101_1_01_001_101_110_0_x_00;
      patterns[2781] = 32'b1010011000010101_1_10_001_101_110_0_x_00;
      patterns[2782] = 32'b1011011000010101_1_11_001_101_110_0_x_00;
      patterns[2783] = 32'b0101011000010000_1_xx_001_xxx_110_0_1_01;
      patterns[2784] = 32'b0100011000010000_0_xx_001_110_xxx_1_x_xx;
      patterns[2785] = 32'b0000011001101001_1_xx_xxx_xxx_110_0_x_10;
      patterns[2786] = 32'b1000011000010110_1_00_001_110_110_0_x_00;
      patterns[2787] = 32'b1001011000010110_1_01_001_110_110_0_x_00;
      patterns[2788] = 32'b1010011000010110_1_10_001_110_110_0_x_00;
      patterns[2789] = 32'b1011011000010110_1_11_001_110_110_0_x_00;
      patterns[2790] = 32'b0101011000010000_1_xx_001_xxx_110_0_1_01;
      patterns[2791] = 32'b0100011000010000_0_xx_001_110_xxx_1_x_xx;
      patterns[2792] = 32'b0000011000110101_1_xx_xxx_xxx_110_0_x_10;
      patterns[2793] = 32'b1000011000010111_1_00_001_111_110_0_x_00;
      patterns[2794] = 32'b1001011000010111_1_01_001_111_110_0_x_00;
      patterns[2795] = 32'b1010011000010111_1_10_001_111_110_0_x_00;
      patterns[2796] = 32'b1011011000010111_1_11_001_111_110_0_x_00;
      patterns[2797] = 32'b0101011000010000_1_xx_001_xxx_110_0_1_01;
      patterns[2798] = 32'b0100011000010000_0_xx_001_110_xxx_1_x_xx;
      patterns[2799] = 32'b0000011001110001_1_xx_xxx_xxx_110_0_x_10;
      patterns[2800] = 32'b1000011000100000_1_00_010_000_110_0_x_00;
      patterns[2801] = 32'b1001011000100000_1_01_010_000_110_0_x_00;
      patterns[2802] = 32'b1010011000100000_1_10_010_000_110_0_x_00;
      patterns[2803] = 32'b1011011000100000_1_11_010_000_110_0_x_00;
      patterns[2804] = 32'b0101011000100000_1_xx_010_xxx_110_0_1_01;
      patterns[2805] = 32'b0100011000100000_0_xx_010_110_xxx_1_x_xx;
      patterns[2806] = 32'b0000011011000101_1_xx_xxx_xxx_110_0_x_10;
      patterns[2807] = 32'b1000011000100001_1_00_010_001_110_0_x_00;
      patterns[2808] = 32'b1001011000100001_1_01_010_001_110_0_x_00;
      patterns[2809] = 32'b1010011000100001_1_10_010_001_110_0_x_00;
      patterns[2810] = 32'b1011011000100001_1_11_010_001_110_0_x_00;
      patterns[2811] = 32'b0101011000100000_1_xx_010_xxx_110_0_1_01;
      patterns[2812] = 32'b0100011000100000_0_xx_010_110_xxx_1_x_xx;
      patterns[2813] = 32'b0000011011111101_1_xx_xxx_xxx_110_0_x_10;
      patterns[2814] = 32'b1000011000100010_1_00_010_010_110_0_x_00;
      patterns[2815] = 32'b1001011000100010_1_01_010_010_110_0_x_00;
      patterns[2816] = 32'b1010011000100010_1_10_010_010_110_0_x_00;
      patterns[2817] = 32'b1011011000100010_1_11_010_010_110_0_x_00;
      patterns[2818] = 32'b0101011000100000_1_xx_010_xxx_110_0_1_01;
      patterns[2819] = 32'b0100011000100000_0_xx_010_110_xxx_1_x_xx;
      patterns[2820] = 32'b0000011000110000_1_xx_xxx_xxx_110_0_x_10;
      patterns[2821] = 32'b1000011000100011_1_00_010_011_110_0_x_00;
      patterns[2822] = 32'b1001011000100011_1_01_010_011_110_0_x_00;
      patterns[2823] = 32'b1010011000100011_1_10_010_011_110_0_x_00;
      patterns[2824] = 32'b1011011000100011_1_11_010_011_110_0_x_00;
      patterns[2825] = 32'b0101011000100000_1_xx_010_xxx_110_0_1_01;
      patterns[2826] = 32'b0100011000100000_0_xx_010_110_xxx_1_x_xx;
      patterns[2827] = 32'b0000011011111110_1_xx_xxx_xxx_110_0_x_10;
      patterns[2828] = 32'b1000011000100100_1_00_010_100_110_0_x_00;
      patterns[2829] = 32'b1001011000100100_1_01_010_100_110_0_x_00;
      patterns[2830] = 32'b1010011000100100_1_10_010_100_110_0_x_00;
      patterns[2831] = 32'b1011011000100100_1_11_010_100_110_0_x_00;
      patterns[2832] = 32'b0101011000100000_1_xx_010_xxx_110_0_1_01;
      patterns[2833] = 32'b0100011000100000_0_xx_010_110_xxx_1_x_xx;
      patterns[2834] = 32'b0000011000110100_1_xx_xxx_xxx_110_0_x_10;
      patterns[2835] = 32'b1000011000100101_1_00_010_101_110_0_x_00;
      patterns[2836] = 32'b1001011000100101_1_01_010_101_110_0_x_00;
      patterns[2837] = 32'b1010011000100101_1_10_010_101_110_0_x_00;
      patterns[2838] = 32'b1011011000100101_1_11_010_101_110_0_x_00;
      patterns[2839] = 32'b0101011000100000_1_xx_010_xxx_110_0_1_01;
      patterns[2840] = 32'b0100011000100000_0_xx_010_110_xxx_1_x_xx;
      patterns[2841] = 32'b0000011010000100_1_xx_xxx_xxx_110_0_x_10;
      patterns[2842] = 32'b1000011000100110_1_00_010_110_110_0_x_00;
      patterns[2843] = 32'b1001011000100110_1_01_010_110_110_0_x_00;
      patterns[2844] = 32'b1010011000100110_1_10_010_110_110_0_x_00;
      patterns[2845] = 32'b1011011000100110_1_11_010_110_110_0_x_00;
      patterns[2846] = 32'b0101011000100000_1_xx_010_xxx_110_0_1_01;
      patterns[2847] = 32'b0100011000100000_0_xx_010_110_xxx_1_x_xx;
      patterns[2848] = 32'b0000011011100111_1_xx_xxx_xxx_110_0_x_10;
      patterns[2849] = 32'b1000011000100111_1_00_010_111_110_0_x_00;
      patterns[2850] = 32'b1001011000100111_1_01_010_111_110_0_x_00;
      patterns[2851] = 32'b1010011000100111_1_10_010_111_110_0_x_00;
      patterns[2852] = 32'b1011011000100111_1_11_010_111_110_0_x_00;
      patterns[2853] = 32'b0101011000100000_1_xx_010_xxx_110_0_1_01;
      patterns[2854] = 32'b0100011000100000_0_xx_010_110_xxx_1_x_xx;
      patterns[2855] = 32'b0000011011110101_1_xx_xxx_xxx_110_0_x_10;
      patterns[2856] = 32'b1000011000110000_1_00_011_000_110_0_x_00;
      patterns[2857] = 32'b1001011000110000_1_01_011_000_110_0_x_00;
      patterns[2858] = 32'b1010011000110000_1_10_011_000_110_0_x_00;
      patterns[2859] = 32'b1011011000110000_1_11_011_000_110_0_x_00;
      patterns[2860] = 32'b0101011000110000_1_xx_011_xxx_110_0_1_01;
      patterns[2861] = 32'b0100011000110000_0_xx_011_110_xxx_1_x_xx;
      patterns[2862] = 32'b0000011001011110_1_xx_xxx_xxx_110_0_x_10;
      patterns[2863] = 32'b1000011000110001_1_00_011_001_110_0_x_00;
      patterns[2864] = 32'b1001011000110001_1_01_011_001_110_0_x_00;
      patterns[2865] = 32'b1010011000110001_1_10_011_001_110_0_x_00;
      patterns[2866] = 32'b1011011000110001_1_11_011_001_110_0_x_00;
      patterns[2867] = 32'b0101011000110000_1_xx_011_xxx_110_0_1_01;
      patterns[2868] = 32'b0100011000110000_0_xx_011_110_xxx_1_x_xx;
      patterns[2869] = 32'b0000011001011100_1_xx_xxx_xxx_110_0_x_10;
      patterns[2870] = 32'b1000011000110010_1_00_011_010_110_0_x_00;
      patterns[2871] = 32'b1001011000110010_1_01_011_010_110_0_x_00;
      patterns[2872] = 32'b1010011000110010_1_10_011_010_110_0_x_00;
      patterns[2873] = 32'b1011011000110010_1_11_011_010_110_0_x_00;
      patterns[2874] = 32'b0101011000110000_1_xx_011_xxx_110_0_1_01;
      patterns[2875] = 32'b0100011000110000_0_xx_011_110_xxx_1_x_xx;
      patterns[2876] = 32'b0000011001110001_1_xx_xxx_xxx_110_0_x_10;
      patterns[2877] = 32'b1000011000110011_1_00_011_011_110_0_x_00;
      patterns[2878] = 32'b1001011000110011_1_01_011_011_110_0_x_00;
      patterns[2879] = 32'b1010011000110011_1_10_011_011_110_0_x_00;
      patterns[2880] = 32'b1011011000110011_1_11_011_011_110_0_x_00;
      patterns[2881] = 32'b0101011000110000_1_xx_011_xxx_110_0_1_01;
      patterns[2882] = 32'b0100011000110000_0_xx_011_110_xxx_1_x_xx;
      patterns[2883] = 32'b0000011011000010_1_xx_xxx_xxx_110_0_x_10;
      patterns[2884] = 32'b1000011000110100_1_00_011_100_110_0_x_00;
      patterns[2885] = 32'b1001011000110100_1_01_011_100_110_0_x_00;
      patterns[2886] = 32'b1010011000110100_1_10_011_100_110_0_x_00;
      patterns[2887] = 32'b1011011000110100_1_11_011_100_110_0_x_00;
      patterns[2888] = 32'b0101011000110000_1_xx_011_xxx_110_0_1_01;
      patterns[2889] = 32'b0100011000110000_0_xx_011_110_xxx_1_x_xx;
      patterns[2890] = 32'b0000011011000101_1_xx_xxx_xxx_110_0_x_10;
      patterns[2891] = 32'b1000011000110101_1_00_011_101_110_0_x_00;
      patterns[2892] = 32'b1001011000110101_1_01_011_101_110_0_x_00;
      patterns[2893] = 32'b1010011000110101_1_10_011_101_110_0_x_00;
      patterns[2894] = 32'b1011011000110101_1_11_011_101_110_0_x_00;
      patterns[2895] = 32'b0101011000110000_1_xx_011_xxx_110_0_1_01;
      patterns[2896] = 32'b0100011000110000_0_xx_011_110_xxx_1_x_xx;
      patterns[2897] = 32'b0000011011010100_1_xx_xxx_xxx_110_0_x_10;
      patterns[2898] = 32'b1000011000110110_1_00_011_110_110_0_x_00;
      patterns[2899] = 32'b1001011000110110_1_01_011_110_110_0_x_00;
      patterns[2900] = 32'b1010011000110110_1_10_011_110_110_0_x_00;
      patterns[2901] = 32'b1011011000110110_1_11_011_110_110_0_x_00;
      patterns[2902] = 32'b0101011000110000_1_xx_011_xxx_110_0_1_01;
      patterns[2903] = 32'b0100011000110000_0_xx_011_110_xxx_1_x_xx;
      patterns[2904] = 32'b0000011001011100_1_xx_xxx_xxx_110_0_x_10;
      patterns[2905] = 32'b1000011000110111_1_00_011_111_110_0_x_00;
      patterns[2906] = 32'b1001011000110111_1_01_011_111_110_0_x_00;
      patterns[2907] = 32'b1010011000110111_1_10_011_111_110_0_x_00;
      patterns[2908] = 32'b1011011000110111_1_11_011_111_110_0_x_00;
      patterns[2909] = 32'b0101011000110000_1_xx_011_xxx_110_0_1_01;
      patterns[2910] = 32'b0100011000110000_0_xx_011_110_xxx_1_x_xx;
      patterns[2911] = 32'b0000011011111110_1_xx_xxx_xxx_110_0_x_10;
      patterns[2912] = 32'b1000011001000000_1_00_100_000_110_0_x_00;
      patterns[2913] = 32'b1001011001000000_1_01_100_000_110_0_x_00;
      patterns[2914] = 32'b1010011001000000_1_10_100_000_110_0_x_00;
      patterns[2915] = 32'b1011011001000000_1_11_100_000_110_0_x_00;
      patterns[2916] = 32'b0101011001000000_1_xx_100_xxx_110_0_1_01;
      patterns[2917] = 32'b0100011001000000_0_xx_100_110_xxx_1_x_xx;
      patterns[2918] = 32'b0000011010000000_1_xx_xxx_xxx_110_0_x_10;
      patterns[2919] = 32'b1000011001000001_1_00_100_001_110_0_x_00;
      patterns[2920] = 32'b1001011001000001_1_01_100_001_110_0_x_00;
      patterns[2921] = 32'b1010011001000001_1_10_100_001_110_0_x_00;
      patterns[2922] = 32'b1011011001000001_1_11_100_001_110_0_x_00;
      patterns[2923] = 32'b0101011001000000_1_xx_100_xxx_110_0_1_01;
      patterns[2924] = 32'b0100011001000000_0_xx_100_110_xxx_1_x_xx;
      patterns[2925] = 32'b0000011000110101_1_xx_xxx_xxx_110_0_x_10;
      patterns[2926] = 32'b1000011001000010_1_00_100_010_110_0_x_00;
      patterns[2927] = 32'b1001011001000010_1_01_100_010_110_0_x_00;
      patterns[2928] = 32'b1010011001000010_1_10_100_010_110_0_x_00;
      patterns[2929] = 32'b1011011001000010_1_11_100_010_110_0_x_00;
      patterns[2930] = 32'b0101011001000000_1_xx_100_xxx_110_0_1_01;
      patterns[2931] = 32'b0100011001000000_0_xx_100_110_xxx_1_x_xx;
      patterns[2932] = 32'b0000011010011010_1_xx_xxx_xxx_110_0_x_10;
      patterns[2933] = 32'b1000011001000011_1_00_100_011_110_0_x_00;
      patterns[2934] = 32'b1001011001000011_1_01_100_011_110_0_x_00;
      patterns[2935] = 32'b1010011001000011_1_10_100_011_110_0_x_00;
      patterns[2936] = 32'b1011011001000011_1_11_100_011_110_0_x_00;
      patterns[2937] = 32'b0101011001000000_1_xx_100_xxx_110_0_1_01;
      patterns[2938] = 32'b0100011001000000_0_xx_100_110_xxx_1_x_xx;
      patterns[2939] = 32'b0000011000101011_1_xx_xxx_xxx_110_0_x_10;
      patterns[2940] = 32'b1000011001000100_1_00_100_100_110_0_x_00;
      patterns[2941] = 32'b1001011001000100_1_01_100_100_110_0_x_00;
      patterns[2942] = 32'b1010011001000100_1_10_100_100_110_0_x_00;
      patterns[2943] = 32'b1011011001000100_1_11_100_100_110_0_x_00;
      patterns[2944] = 32'b0101011001000000_1_xx_100_xxx_110_0_1_01;
      patterns[2945] = 32'b0100011001000000_0_xx_100_110_xxx_1_x_xx;
      patterns[2946] = 32'b0000011011000100_1_xx_xxx_xxx_110_0_x_10;
      patterns[2947] = 32'b1000011001000101_1_00_100_101_110_0_x_00;
      patterns[2948] = 32'b1001011001000101_1_01_100_101_110_0_x_00;
      patterns[2949] = 32'b1010011001000101_1_10_100_101_110_0_x_00;
      patterns[2950] = 32'b1011011001000101_1_11_100_101_110_0_x_00;
      patterns[2951] = 32'b0101011001000000_1_xx_100_xxx_110_0_1_01;
      patterns[2952] = 32'b0100011001000000_0_xx_100_110_xxx_1_x_xx;
      patterns[2953] = 32'b0000011010100010_1_xx_xxx_xxx_110_0_x_10;
      patterns[2954] = 32'b1000011001000110_1_00_100_110_110_0_x_00;
      patterns[2955] = 32'b1001011001000110_1_01_100_110_110_0_x_00;
      patterns[2956] = 32'b1010011001000110_1_10_100_110_110_0_x_00;
      patterns[2957] = 32'b1011011001000110_1_11_100_110_110_0_x_00;
      patterns[2958] = 32'b0101011001000000_1_xx_100_xxx_110_0_1_01;
      patterns[2959] = 32'b0100011001000000_0_xx_100_110_xxx_1_x_xx;
      patterns[2960] = 32'b0000011001011101_1_xx_xxx_xxx_110_0_x_10;
      patterns[2961] = 32'b1000011001000111_1_00_100_111_110_0_x_00;
      patterns[2962] = 32'b1001011001000111_1_01_100_111_110_0_x_00;
      patterns[2963] = 32'b1010011001000111_1_10_100_111_110_0_x_00;
      patterns[2964] = 32'b1011011001000111_1_11_100_111_110_0_x_00;
      patterns[2965] = 32'b0101011001000000_1_xx_100_xxx_110_0_1_01;
      patterns[2966] = 32'b0100011001000000_0_xx_100_110_xxx_1_x_xx;
      patterns[2967] = 32'b0000011000010110_1_xx_xxx_xxx_110_0_x_10;
      patterns[2968] = 32'b1000011001010000_1_00_101_000_110_0_x_00;
      patterns[2969] = 32'b1001011001010000_1_01_101_000_110_0_x_00;
      patterns[2970] = 32'b1010011001010000_1_10_101_000_110_0_x_00;
      patterns[2971] = 32'b1011011001010000_1_11_101_000_110_0_x_00;
      patterns[2972] = 32'b0101011001010000_1_xx_101_xxx_110_0_1_01;
      patterns[2973] = 32'b0100011001010000_0_xx_101_110_xxx_1_x_xx;
      patterns[2974] = 32'b0000011001101010_1_xx_xxx_xxx_110_0_x_10;
      patterns[2975] = 32'b1000011001010001_1_00_101_001_110_0_x_00;
      patterns[2976] = 32'b1001011001010001_1_01_101_001_110_0_x_00;
      patterns[2977] = 32'b1010011001010001_1_10_101_001_110_0_x_00;
      patterns[2978] = 32'b1011011001010001_1_11_101_001_110_0_x_00;
      patterns[2979] = 32'b0101011001010000_1_xx_101_xxx_110_0_1_01;
      patterns[2980] = 32'b0100011001010000_0_xx_101_110_xxx_1_x_xx;
      patterns[2981] = 32'b0000011001001000_1_xx_xxx_xxx_110_0_x_10;
      patterns[2982] = 32'b1000011001010010_1_00_101_010_110_0_x_00;
      patterns[2983] = 32'b1001011001010010_1_01_101_010_110_0_x_00;
      patterns[2984] = 32'b1010011001010010_1_10_101_010_110_0_x_00;
      patterns[2985] = 32'b1011011001010010_1_11_101_010_110_0_x_00;
      patterns[2986] = 32'b0101011001010000_1_xx_101_xxx_110_0_1_01;
      patterns[2987] = 32'b0100011001010000_0_xx_101_110_xxx_1_x_xx;
      patterns[2988] = 32'b0000011010100011_1_xx_xxx_xxx_110_0_x_10;
      patterns[2989] = 32'b1000011001010011_1_00_101_011_110_0_x_00;
      patterns[2990] = 32'b1001011001010011_1_01_101_011_110_0_x_00;
      patterns[2991] = 32'b1010011001010011_1_10_101_011_110_0_x_00;
      patterns[2992] = 32'b1011011001010011_1_11_101_011_110_0_x_00;
      patterns[2993] = 32'b0101011001010000_1_xx_101_xxx_110_0_1_01;
      patterns[2994] = 32'b0100011001010000_0_xx_101_110_xxx_1_x_xx;
      patterns[2995] = 32'b0000011010110101_1_xx_xxx_xxx_110_0_x_10;
      patterns[2996] = 32'b1000011001010100_1_00_101_100_110_0_x_00;
      patterns[2997] = 32'b1001011001010100_1_01_101_100_110_0_x_00;
      patterns[2998] = 32'b1010011001010100_1_10_101_100_110_0_x_00;
      patterns[2999] = 32'b1011011001010100_1_11_101_100_110_0_x_00;
      patterns[3000] = 32'b0101011001010000_1_xx_101_xxx_110_0_1_01;
      patterns[3001] = 32'b0100011001010000_0_xx_101_110_xxx_1_x_xx;
      patterns[3002] = 32'b0000011001001100_1_xx_xxx_xxx_110_0_x_10;
      patterns[3003] = 32'b1000011001010101_1_00_101_101_110_0_x_00;
      patterns[3004] = 32'b1001011001010101_1_01_101_101_110_0_x_00;
      patterns[3005] = 32'b1010011001010101_1_10_101_101_110_0_x_00;
      patterns[3006] = 32'b1011011001010101_1_11_101_101_110_0_x_00;
      patterns[3007] = 32'b0101011001010000_1_xx_101_xxx_110_0_1_01;
      patterns[3008] = 32'b0100011001010000_0_xx_101_110_xxx_1_x_xx;
      patterns[3009] = 32'b0000011000111000_1_xx_xxx_xxx_110_0_x_10;
      patterns[3010] = 32'b1000011001010110_1_00_101_110_110_0_x_00;
      patterns[3011] = 32'b1001011001010110_1_01_101_110_110_0_x_00;
      patterns[3012] = 32'b1010011001010110_1_10_101_110_110_0_x_00;
      patterns[3013] = 32'b1011011001010110_1_11_101_110_110_0_x_00;
      patterns[3014] = 32'b0101011001010000_1_xx_101_xxx_110_0_1_01;
      patterns[3015] = 32'b0100011001010000_0_xx_101_110_xxx_1_x_xx;
      patterns[3016] = 32'b0000011011101001_1_xx_xxx_xxx_110_0_x_10;
      patterns[3017] = 32'b1000011001010111_1_00_101_111_110_0_x_00;
      patterns[3018] = 32'b1001011001010111_1_01_101_111_110_0_x_00;
      patterns[3019] = 32'b1010011001010111_1_10_101_111_110_0_x_00;
      patterns[3020] = 32'b1011011001010111_1_11_101_111_110_0_x_00;
      patterns[3021] = 32'b0101011001010000_1_xx_101_xxx_110_0_1_01;
      patterns[3022] = 32'b0100011001010000_0_xx_101_110_xxx_1_x_xx;
      patterns[3023] = 32'b0000011011100000_1_xx_xxx_xxx_110_0_x_10;
      patterns[3024] = 32'b1000011001100000_1_00_110_000_110_0_x_00;
      patterns[3025] = 32'b1001011001100000_1_01_110_000_110_0_x_00;
      patterns[3026] = 32'b1010011001100000_1_10_110_000_110_0_x_00;
      patterns[3027] = 32'b1011011001100000_1_11_110_000_110_0_x_00;
      patterns[3028] = 32'b0101011001100000_1_xx_110_xxx_110_0_1_01;
      patterns[3029] = 32'b0100011001100000_0_xx_110_110_xxx_1_x_xx;
      patterns[3030] = 32'b0000011000000100_1_xx_xxx_xxx_110_0_x_10;
      patterns[3031] = 32'b1000011001100001_1_00_110_001_110_0_x_00;
      patterns[3032] = 32'b1001011001100001_1_01_110_001_110_0_x_00;
      patterns[3033] = 32'b1010011001100001_1_10_110_001_110_0_x_00;
      patterns[3034] = 32'b1011011001100001_1_11_110_001_110_0_x_00;
      patterns[3035] = 32'b0101011001100000_1_xx_110_xxx_110_0_1_01;
      patterns[3036] = 32'b0100011001100000_0_xx_110_110_xxx_1_x_xx;
      patterns[3037] = 32'b0000011000000000_1_xx_xxx_xxx_110_0_x_10;
      patterns[3038] = 32'b1000011001100010_1_00_110_010_110_0_x_00;
      patterns[3039] = 32'b1001011001100010_1_01_110_010_110_0_x_00;
      patterns[3040] = 32'b1010011001100010_1_10_110_010_110_0_x_00;
      patterns[3041] = 32'b1011011001100010_1_11_110_010_110_0_x_00;
      patterns[3042] = 32'b0101011001100000_1_xx_110_xxx_110_0_1_01;
      patterns[3043] = 32'b0100011001100000_0_xx_110_110_xxx_1_x_xx;
      patterns[3044] = 32'b0000011011100000_1_xx_xxx_xxx_110_0_x_10;
      patterns[3045] = 32'b1000011001100011_1_00_110_011_110_0_x_00;
      patterns[3046] = 32'b1001011001100011_1_01_110_011_110_0_x_00;
      patterns[3047] = 32'b1010011001100011_1_10_110_011_110_0_x_00;
      patterns[3048] = 32'b1011011001100011_1_11_110_011_110_0_x_00;
      patterns[3049] = 32'b0101011001100000_1_xx_110_xxx_110_0_1_01;
      patterns[3050] = 32'b0100011001100000_0_xx_110_110_xxx_1_x_xx;
      patterns[3051] = 32'b0000011000000100_1_xx_xxx_xxx_110_0_x_10;
      patterns[3052] = 32'b1000011001100100_1_00_110_100_110_0_x_00;
      patterns[3053] = 32'b1001011001100100_1_01_110_100_110_0_x_00;
      patterns[3054] = 32'b1010011001100100_1_10_110_100_110_0_x_00;
      patterns[3055] = 32'b1011011001100100_1_11_110_100_110_0_x_00;
      patterns[3056] = 32'b0101011001100000_1_xx_110_xxx_110_0_1_01;
      patterns[3057] = 32'b0100011001100000_0_xx_110_110_xxx_1_x_xx;
      patterns[3058] = 32'b0000011011011000_1_xx_xxx_xxx_110_0_x_10;
      patterns[3059] = 32'b1000011001100101_1_00_110_101_110_0_x_00;
      patterns[3060] = 32'b1001011001100101_1_01_110_101_110_0_x_00;
      patterns[3061] = 32'b1010011001100101_1_10_110_101_110_0_x_00;
      patterns[3062] = 32'b1011011001100101_1_11_110_101_110_0_x_00;
      patterns[3063] = 32'b0101011001100000_1_xx_110_xxx_110_0_1_01;
      patterns[3064] = 32'b0100011001100000_0_xx_110_110_xxx_1_x_xx;
      patterns[3065] = 32'b0000011010100011_1_xx_xxx_xxx_110_0_x_10;
      patterns[3066] = 32'b1000011001100110_1_00_110_110_110_0_x_00;
      patterns[3067] = 32'b1001011001100110_1_01_110_110_110_0_x_00;
      patterns[3068] = 32'b1010011001100110_1_10_110_110_110_0_x_00;
      patterns[3069] = 32'b1011011001100110_1_11_110_110_110_0_x_00;
      patterns[3070] = 32'b0101011001100000_1_xx_110_xxx_110_0_1_01;
      patterns[3071] = 32'b0100011001100000_0_xx_110_110_xxx_1_x_xx;
      patterns[3072] = 32'b0000011000001000_1_xx_xxx_xxx_110_0_x_10;
      patterns[3073] = 32'b1000011001100111_1_00_110_111_110_0_x_00;
      patterns[3074] = 32'b1001011001100111_1_01_110_111_110_0_x_00;
      patterns[3075] = 32'b1010011001100111_1_10_110_111_110_0_x_00;
      patterns[3076] = 32'b1011011001100111_1_11_110_111_110_0_x_00;
      patterns[3077] = 32'b0101011001100000_1_xx_110_xxx_110_0_1_01;
      patterns[3078] = 32'b0100011001100000_0_xx_110_110_xxx_1_x_xx;
      patterns[3079] = 32'b0000011000111011_1_xx_xxx_xxx_110_0_x_10;
      patterns[3080] = 32'b1000011001110000_1_00_111_000_110_0_x_00;
      patterns[3081] = 32'b1001011001110000_1_01_111_000_110_0_x_00;
      patterns[3082] = 32'b1010011001110000_1_10_111_000_110_0_x_00;
      patterns[3083] = 32'b1011011001110000_1_11_111_000_110_0_x_00;
      patterns[3084] = 32'b0101011001110000_1_xx_111_xxx_110_0_1_01;
      patterns[3085] = 32'b0100011001110000_0_xx_111_110_xxx_1_x_xx;
      patterns[3086] = 32'b0000011011000010_1_xx_xxx_xxx_110_0_x_10;
      patterns[3087] = 32'b1000011001110001_1_00_111_001_110_0_x_00;
      patterns[3088] = 32'b1001011001110001_1_01_111_001_110_0_x_00;
      patterns[3089] = 32'b1010011001110001_1_10_111_001_110_0_x_00;
      patterns[3090] = 32'b1011011001110001_1_11_111_001_110_0_x_00;
      patterns[3091] = 32'b0101011001110000_1_xx_111_xxx_110_0_1_01;
      patterns[3092] = 32'b0100011001110000_0_xx_111_110_xxx_1_x_xx;
      patterns[3093] = 32'b0000011001010111_1_xx_xxx_xxx_110_0_x_10;
      patterns[3094] = 32'b1000011001110010_1_00_111_010_110_0_x_00;
      patterns[3095] = 32'b1001011001110010_1_01_111_010_110_0_x_00;
      patterns[3096] = 32'b1010011001110010_1_10_111_010_110_0_x_00;
      patterns[3097] = 32'b1011011001110010_1_11_111_010_110_0_x_00;
      patterns[3098] = 32'b0101011001110000_1_xx_111_xxx_110_0_1_01;
      patterns[3099] = 32'b0100011001110000_0_xx_111_110_xxx_1_x_xx;
      patterns[3100] = 32'b0000011011000100_1_xx_xxx_xxx_110_0_x_10;
      patterns[3101] = 32'b1000011001110011_1_00_111_011_110_0_x_00;
      patterns[3102] = 32'b1001011001110011_1_01_111_011_110_0_x_00;
      patterns[3103] = 32'b1010011001110011_1_10_111_011_110_0_x_00;
      patterns[3104] = 32'b1011011001110011_1_11_111_011_110_0_x_00;
      patterns[3105] = 32'b0101011001110000_1_xx_111_xxx_110_0_1_01;
      patterns[3106] = 32'b0100011001110000_0_xx_111_110_xxx_1_x_xx;
      patterns[3107] = 32'b0000011010111110_1_xx_xxx_xxx_110_0_x_10;
      patterns[3108] = 32'b1000011001110100_1_00_111_100_110_0_x_00;
      patterns[3109] = 32'b1001011001110100_1_01_111_100_110_0_x_00;
      patterns[3110] = 32'b1010011001110100_1_10_111_100_110_0_x_00;
      patterns[3111] = 32'b1011011001110100_1_11_111_100_110_0_x_00;
      patterns[3112] = 32'b0101011001110000_1_xx_111_xxx_110_0_1_01;
      patterns[3113] = 32'b0100011001110000_0_xx_111_110_xxx_1_x_xx;
      patterns[3114] = 32'b0000011011101000_1_xx_xxx_xxx_110_0_x_10;
      patterns[3115] = 32'b1000011001110101_1_00_111_101_110_0_x_00;
      patterns[3116] = 32'b1001011001110101_1_01_111_101_110_0_x_00;
      patterns[3117] = 32'b1010011001110101_1_10_111_101_110_0_x_00;
      patterns[3118] = 32'b1011011001110101_1_11_111_101_110_0_x_00;
      patterns[3119] = 32'b0101011001110000_1_xx_111_xxx_110_0_1_01;
      patterns[3120] = 32'b0100011001110000_0_xx_111_110_xxx_1_x_xx;
      patterns[3121] = 32'b0000011010011101_1_xx_xxx_xxx_110_0_x_10;
      patterns[3122] = 32'b1000011001110110_1_00_111_110_110_0_x_00;
      patterns[3123] = 32'b1001011001110110_1_01_111_110_110_0_x_00;
      patterns[3124] = 32'b1010011001110110_1_10_111_110_110_0_x_00;
      patterns[3125] = 32'b1011011001110110_1_11_111_110_110_0_x_00;
      patterns[3126] = 32'b0101011001110000_1_xx_111_xxx_110_0_1_01;
      patterns[3127] = 32'b0100011001110000_0_xx_111_110_xxx_1_x_xx;
      patterns[3128] = 32'b0000011011001110_1_xx_xxx_xxx_110_0_x_10;
      patterns[3129] = 32'b1000011001110111_1_00_111_111_110_0_x_00;
      patterns[3130] = 32'b1001011001110111_1_01_111_111_110_0_x_00;
      patterns[3131] = 32'b1010011001110111_1_10_111_111_110_0_x_00;
      patterns[3132] = 32'b1011011001110111_1_11_111_111_110_0_x_00;
      patterns[3133] = 32'b0101011001110000_1_xx_111_xxx_110_0_1_01;
      patterns[3134] = 32'b0100011001110000_0_xx_111_110_xxx_1_x_xx;
      patterns[3135] = 32'b0000011011001001_1_xx_xxx_xxx_110_0_x_10;
      patterns[3136] = 32'b1000011100000000_1_00_000_000_111_0_x_00;
      patterns[3137] = 32'b1001011100000000_1_01_000_000_111_0_x_00;
      patterns[3138] = 32'b1010011100000000_1_10_000_000_111_0_x_00;
      patterns[3139] = 32'b1011011100000000_1_11_000_000_111_0_x_00;
      patterns[3140] = 32'b0101011100000000_1_xx_000_xxx_111_0_1_01;
      patterns[3141] = 32'b0100011100000000_0_xx_000_111_xxx_1_x_xx;
      patterns[3142] = 32'b0000011101101110_1_xx_xxx_xxx_111_0_x_10;
      patterns[3143] = 32'b1000011100000001_1_00_000_001_111_0_x_00;
      patterns[3144] = 32'b1001011100000001_1_01_000_001_111_0_x_00;
      patterns[3145] = 32'b1010011100000001_1_10_000_001_111_0_x_00;
      patterns[3146] = 32'b1011011100000001_1_11_000_001_111_0_x_00;
      patterns[3147] = 32'b0101011100000000_1_xx_000_xxx_111_0_1_01;
      patterns[3148] = 32'b0100011100000000_0_xx_000_111_xxx_1_x_xx;
      patterns[3149] = 32'b0000011111101000_1_xx_xxx_xxx_111_0_x_10;
      patterns[3150] = 32'b1000011100000010_1_00_000_010_111_0_x_00;
      patterns[3151] = 32'b1001011100000010_1_01_000_010_111_0_x_00;
      patterns[3152] = 32'b1010011100000010_1_10_000_010_111_0_x_00;
      patterns[3153] = 32'b1011011100000010_1_11_000_010_111_0_x_00;
      patterns[3154] = 32'b0101011100000000_1_xx_000_xxx_111_0_1_01;
      patterns[3155] = 32'b0100011100000000_0_xx_000_111_xxx_1_x_xx;
      patterns[3156] = 32'b0000011111100110_1_xx_xxx_xxx_111_0_x_10;
      patterns[3157] = 32'b1000011100000011_1_00_000_011_111_0_x_00;
      patterns[3158] = 32'b1001011100000011_1_01_000_011_111_0_x_00;
      patterns[3159] = 32'b1010011100000011_1_10_000_011_111_0_x_00;
      patterns[3160] = 32'b1011011100000011_1_11_000_011_111_0_x_00;
      patterns[3161] = 32'b0101011100000000_1_xx_000_xxx_111_0_1_01;
      patterns[3162] = 32'b0100011100000000_0_xx_000_111_xxx_1_x_xx;
      patterns[3163] = 32'b0000011101010111_1_xx_xxx_xxx_111_0_x_10;
      patterns[3164] = 32'b1000011100000100_1_00_000_100_111_0_x_00;
      patterns[3165] = 32'b1001011100000100_1_01_000_100_111_0_x_00;
      patterns[3166] = 32'b1010011100000100_1_10_000_100_111_0_x_00;
      patterns[3167] = 32'b1011011100000100_1_11_000_100_111_0_x_00;
      patterns[3168] = 32'b0101011100000000_1_xx_000_xxx_111_0_1_01;
      patterns[3169] = 32'b0100011100000000_0_xx_000_111_xxx_1_x_xx;
      patterns[3170] = 32'b0000011100101101_1_xx_xxx_xxx_111_0_x_10;
      patterns[3171] = 32'b1000011100000101_1_00_000_101_111_0_x_00;
      patterns[3172] = 32'b1001011100000101_1_01_000_101_111_0_x_00;
      patterns[3173] = 32'b1010011100000101_1_10_000_101_111_0_x_00;
      patterns[3174] = 32'b1011011100000101_1_11_000_101_111_0_x_00;
      patterns[3175] = 32'b0101011100000000_1_xx_000_xxx_111_0_1_01;
      patterns[3176] = 32'b0100011100000000_0_xx_000_111_xxx_1_x_xx;
      patterns[3177] = 32'b0000011100010110_1_xx_xxx_xxx_111_0_x_10;
      patterns[3178] = 32'b1000011100000110_1_00_000_110_111_0_x_00;
      patterns[3179] = 32'b1001011100000110_1_01_000_110_111_0_x_00;
      patterns[3180] = 32'b1010011100000110_1_10_000_110_111_0_x_00;
      patterns[3181] = 32'b1011011100000110_1_11_000_110_111_0_x_00;
      patterns[3182] = 32'b0101011100000000_1_xx_000_xxx_111_0_1_01;
      patterns[3183] = 32'b0100011100000000_0_xx_000_111_xxx_1_x_xx;
      patterns[3184] = 32'b0000011101101001_1_xx_xxx_xxx_111_0_x_10;
      patterns[3185] = 32'b1000011100000111_1_00_000_111_111_0_x_00;
      patterns[3186] = 32'b1001011100000111_1_01_000_111_111_0_x_00;
      patterns[3187] = 32'b1010011100000111_1_10_000_111_111_0_x_00;
      patterns[3188] = 32'b1011011100000111_1_11_000_111_111_0_x_00;
      patterns[3189] = 32'b0101011100000000_1_xx_000_xxx_111_0_1_01;
      patterns[3190] = 32'b0100011100000000_0_xx_000_111_xxx_1_x_xx;
      patterns[3191] = 32'b0000011100101000_1_xx_xxx_xxx_111_0_x_10;
      patterns[3192] = 32'b1000011100010000_1_00_001_000_111_0_x_00;
      patterns[3193] = 32'b1001011100010000_1_01_001_000_111_0_x_00;
      patterns[3194] = 32'b1010011100010000_1_10_001_000_111_0_x_00;
      patterns[3195] = 32'b1011011100010000_1_11_001_000_111_0_x_00;
      patterns[3196] = 32'b0101011100010000_1_xx_001_xxx_111_0_1_01;
      patterns[3197] = 32'b0100011100010000_0_xx_001_111_xxx_1_x_xx;
      patterns[3198] = 32'b0000011111010110_1_xx_xxx_xxx_111_0_x_10;
      patterns[3199] = 32'b1000011100010001_1_00_001_001_111_0_x_00;
      patterns[3200] = 32'b1001011100010001_1_01_001_001_111_0_x_00;
      patterns[3201] = 32'b1010011100010001_1_10_001_001_111_0_x_00;
      patterns[3202] = 32'b1011011100010001_1_11_001_001_111_0_x_00;
      patterns[3203] = 32'b0101011100010000_1_xx_001_xxx_111_0_1_01;
      patterns[3204] = 32'b0100011100010000_0_xx_001_111_xxx_1_x_xx;
      patterns[3205] = 32'b0000011101010100_1_xx_xxx_xxx_111_0_x_10;
      patterns[3206] = 32'b1000011100010010_1_00_001_010_111_0_x_00;
      patterns[3207] = 32'b1001011100010010_1_01_001_010_111_0_x_00;
      patterns[3208] = 32'b1010011100010010_1_10_001_010_111_0_x_00;
      patterns[3209] = 32'b1011011100010010_1_11_001_010_111_0_x_00;
      patterns[3210] = 32'b0101011100010000_1_xx_001_xxx_111_0_1_01;
      patterns[3211] = 32'b0100011100010000_0_xx_001_111_xxx_1_x_xx;
      patterns[3212] = 32'b0000011110001001_1_xx_xxx_xxx_111_0_x_10;
      patterns[3213] = 32'b1000011100010011_1_00_001_011_111_0_x_00;
      patterns[3214] = 32'b1001011100010011_1_01_001_011_111_0_x_00;
      patterns[3215] = 32'b1010011100010011_1_10_001_011_111_0_x_00;
      patterns[3216] = 32'b1011011100010011_1_11_001_011_111_0_x_00;
      patterns[3217] = 32'b0101011100010000_1_xx_001_xxx_111_0_1_01;
      patterns[3218] = 32'b0100011100010000_0_xx_001_111_xxx_1_x_xx;
      patterns[3219] = 32'b0000011110001001_1_xx_xxx_xxx_111_0_x_10;
      patterns[3220] = 32'b1000011100010100_1_00_001_100_111_0_x_00;
      patterns[3221] = 32'b1001011100010100_1_01_001_100_111_0_x_00;
      patterns[3222] = 32'b1010011100010100_1_10_001_100_111_0_x_00;
      patterns[3223] = 32'b1011011100010100_1_11_001_100_111_0_x_00;
      patterns[3224] = 32'b0101011100010000_1_xx_001_xxx_111_0_1_01;
      patterns[3225] = 32'b0100011100010000_0_xx_001_111_xxx_1_x_xx;
      patterns[3226] = 32'b0000011111010100_1_xx_xxx_xxx_111_0_x_10;
      patterns[3227] = 32'b1000011100010101_1_00_001_101_111_0_x_00;
      patterns[3228] = 32'b1001011100010101_1_01_001_101_111_0_x_00;
      patterns[3229] = 32'b1010011100010101_1_10_001_101_111_0_x_00;
      patterns[3230] = 32'b1011011100010101_1_11_001_101_111_0_x_00;
      patterns[3231] = 32'b0101011100010000_1_xx_001_xxx_111_0_1_01;
      patterns[3232] = 32'b0100011100010000_0_xx_001_111_xxx_1_x_xx;
      patterns[3233] = 32'b0000011100000000_1_xx_xxx_xxx_111_0_x_10;
      patterns[3234] = 32'b1000011100010110_1_00_001_110_111_0_x_00;
      patterns[3235] = 32'b1001011100010110_1_01_001_110_111_0_x_00;
      patterns[3236] = 32'b1010011100010110_1_10_001_110_111_0_x_00;
      patterns[3237] = 32'b1011011100010110_1_11_001_110_111_0_x_00;
      patterns[3238] = 32'b0101011100010000_1_xx_001_xxx_111_0_1_01;
      patterns[3239] = 32'b0100011100010000_0_xx_001_111_xxx_1_x_xx;
      patterns[3240] = 32'b0000011100011000_1_xx_xxx_xxx_111_0_x_10;
      patterns[3241] = 32'b1000011100010111_1_00_001_111_111_0_x_00;
      patterns[3242] = 32'b1001011100010111_1_01_001_111_111_0_x_00;
      patterns[3243] = 32'b1010011100010111_1_10_001_111_111_0_x_00;
      patterns[3244] = 32'b1011011100010111_1_11_001_111_111_0_x_00;
      patterns[3245] = 32'b0101011100010000_1_xx_001_xxx_111_0_1_01;
      patterns[3246] = 32'b0100011100010000_0_xx_001_111_xxx_1_x_xx;
      patterns[3247] = 32'b0000011100111101_1_xx_xxx_xxx_111_0_x_10;
      patterns[3248] = 32'b1000011100100000_1_00_010_000_111_0_x_00;
      patterns[3249] = 32'b1001011100100000_1_01_010_000_111_0_x_00;
      patterns[3250] = 32'b1010011100100000_1_10_010_000_111_0_x_00;
      patterns[3251] = 32'b1011011100100000_1_11_010_000_111_0_x_00;
      patterns[3252] = 32'b0101011100100000_1_xx_010_xxx_111_0_1_01;
      patterns[3253] = 32'b0100011100100000_0_xx_010_111_xxx_1_x_xx;
      patterns[3254] = 32'b0000011110110001_1_xx_xxx_xxx_111_0_x_10;
      patterns[3255] = 32'b1000011100100001_1_00_010_001_111_0_x_00;
      patterns[3256] = 32'b1001011100100001_1_01_010_001_111_0_x_00;
      patterns[3257] = 32'b1010011100100001_1_10_010_001_111_0_x_00;
      patterns[3258] = 32'b1011011100100001_1_11_010_001_111_0_x_00;
      patterns[3259] = 32'b0101011100100000_1_xx_010_xxx_111_0_1_01;
      patterns[3260] = 32'b0100011100100000_0_xx_010_111_xxx_1_x_xx;
      patterns[3261] = 32'b0000011100110010_1_xx_xxx_xxx_111_0_x_10;
      patterns[3262] = 32'b1000011100100010_1_00_010_010_111_0_x_00;
      patterns[3263] = 32'b1001011100100010_1_01_010_010_111_0_x_00;
      patterns[3264] = 32'b1010011100100010_1_10_010_010_111_0_x_00;
      patterns[3265] = 32'b1011011100100010_1_11_010_010_111_0_x_00;
      patterns[3266] = 32'b0101011100100000_1_xx_010_xxx_111_0_1_01;
      patterns[3267] = 32'b0100011100100000_0_xx_010_111_xxx_1_x_xx;
      patterns[3268] = 32'b0000011101001100_1_xx_xxx_xxx_111_0_x_10;
      patterns[3269] = 32'b1000011100100011_1_00_010_011_111_0_x_00;
      patterns[3270] = 32'b1001011100100011_1_01_010_011_111_0_x_00;
      patterns[3271] = 32'b1010011100100011_1_10_010_011_111_0_x_00;
      patterns[3272] = 32'b1011011100100011_1_11_010_011_111_0_x_00;
      patterns[3273] = 32'b0101011100100000_1_xx_010_xxx_111_0_1_01;
      patterns[3274] = 32'b0100011100100000_0_xx_010_111_xxx_1_x_xx;
      patterns[3275] = 32'b0000011110110011_1_xx_xxx_xxx_111_0_x_10;
      patterns[3276] = 32'b1000011100100100_1_00_010_100_111_0_x_00;
      patterns[3277] = 32'b1001011100100100_1_01_010_100_111_0_x_00;
      patterns[3278] = 32'b1010011100100100_1_10_010_100_111_0_x_00;
      patterns[3279] = 32'b1011011100100100_1_11_010_100_111_0_x_00;
      patterns[3280] = 32'b0101011100100000_1_xx_010_xxx_111_0_1_01;
      patterns[3281] = 32'b0100011100100000_0_xx_010_111_xxx_1_x_xx;
      patterns[3282] = 32'b0000011111011001_1_xx_xxx_xxx_111_0_x_10;
      patterns[3283] = 32'b1000011100100101_1_00_010_101_111_0_x_00;
      patterns[3284] = 32'b1001011100100101_1_01_010_101_111_0_x_00;
      patterns[3285] = 32'b1010011100100101_1_10_010_101_111_0_x_00;
      patterns[3286] = 32'b1011011100100101_1_11_010_101_111_0_x_00;
      patterns[3287] = 32'b0101011100100000_1_xx_010_xxx_111_0_1_01;
      patterns[3288] = 32'b0100011100100000_0_xx_010_111_xxx_1_x_xx;
      patterns[3289] = 32'b0000011101010011_1_xx_xxx_xxx_111_0_x_10;
      patterns[3290] = 32'b1000011100100110_1_00_010_110_111_0_x_00;
      patterns[3291] = 32'b1001011100100110_1_01_010_110_111_0_x_00;
      patterns[3292] = 32'b1010011100100110_1_10_010_110_111_0_x_00;
      patterns[3293] = 32'b1011011100100110_1_11_010_110_111_0_x_00;
      patterns[3294] = 32'b0101011100100000_1_xx_010_xxx_111_0_1_01;
      patterns[3295] = 32'b0100011100100000_0_xx_010_111_xxx_1_x_xx;
      patterns[3296] = 32'b0000011100111111_1_xx_xxx_xxx_111_0_x_10;
      patterns[3297] = 32'b1000011100100111_1_00_010_111_111_0_x_00;
      patterns[3298] = 32'b1001011100100111_1_01_010_111_111_0_x_00;
      patterns[3299] = 32'b1010011100100111_1_10_010_111_111_0_x_00;
      patterns[3300] = 32'b1011011100100111_1_11_010_111_111_0_x_00;
      patterns[3301] = 32'b0101011100100000_1_xx_010_xxx_111_0_1_01;
      patterns[3302] = 32'b0100011100100000_0_xx_010_111_xxx_1_x_xx;
      patterns[3303] = 32'b0000011101110111_1_xx_xxx_xxx_111_0_x_10;
      patterns[3304] = 32'b1000011100110000_1_00_011_000_111_0_x_00;
      patterns[3305] = 32'b1001011100110000_1_01_011_000_111_0_x_00;
      patterns[3306] = 32'b1010011100110000_1_10_011_000_111_0_x_00;
      patterns[3307] = 32'b1011011100110000_1_11_011_000_111_0_x_00;
      patterns[3308] = 32'b0101011100110000_1_xx_011_xxx_111_0_1_01;
      patterns[3309] = 32'b0100011100110000_0_xx_011_111_xxx_1_x_xx;
      patterns[3310] = 32'b0000011100110000_1_xx_xxx_xxx_111_0_x_10;
      patterns[3311] = 32'b1000011100110001_1_00_011_001_111_0_x_00;
      patterns[3312] = 32'b1001011100110001_1_01_011_001_111_0_x_00;
      patterns[3313] = 32'b1010011100110001_1_10_011_001_111_0_x_00;
      patterns[3314] = 32'b1011011100110001_1_11_011_001_111_0_x_00;
      patterns[3315] = 32'b0101011100110000_1_xx_011_xxx_111_0_1_01;
      patterns[3316] = 32'b0100011100110000_0_xx_011_111_xxx_1_x_xx;
      patterns[3317] = 32'b0000011100110001_1_xx_xxx_xxx_111_0_x_10;
      patterns[3318] = 32'b1000011100110010_1_00_011_010_111_0_x_00;
      patterns[3319] = 32'b1001011100110010_1_01_011_010_111_0_x_00;
      patterns[3320] = 32'b1010011100110010_1_10_011_010_111_0_x_00;
      patterns[3321] = 32'b1011011100110010_1_11_011_010_111_0_x_00;
      patterns[3322] = 32'b0101011100110000_1_xx_011_xxx_111_0_1_01;
      patterns[3323] = 32'b0100011100110000_0_xx_011_111_xxx_1_x_xx;
      patterns[3324] = 32'b0000011111001111_1_xx_xxx_xxx_111_0_x_10;
      patterns[3325] = 32'b1000011100110011_1_00_011_011_111_0_x_00;
      patterns[3326] = 32'b1001011100110011_1_01_011_011_111_0_x_00;
      patterns[3327] = 32'b1010011100110011_1_10_011_011_111_0_x_00;
      patterns[3328] = 32'b1011011100110011_1_11_011_011_111_0_x_00;
      patterns[3329] = 32'b0101011100110000_1_xx_011_xxx_111_0_1_01;
      patterns[3330] = 32'b0100011100110000_0_xx_011_111_xxx_1_x_xx;
      patterns[3331] = 32'b0000011101101100_1_xx_xxx_xxx_111_0_x_10;
      patterns[3332] = 32'b1000011100110100_1_00_011_100_111_0_x_00;
      patterns[3333] = 32'b1001011100110100_1_01_011_100_111_0_x_00;
      patterns[3334] = 32'b1010011100110100_1_10_011_100_111_0_x_00;
      patterns[3335] = 32'b1011011100110100_1_11_011_100_111_0_x_00;
      patterns[3336] = 32'b0101011100110000_1_xx_011_xxx_111_0_1_01;
      patterns[3337] = 32'b0100011100110000_0_xx_011_111_xxx_1_x_xx;
      patterns[3338] = 32'b0000011110010000_1_xx_xxx_xxx_111_0_x_10;
      patterns[3339] = 32'b1000011100110101_1_00_011_101_111_0_x_00;
      patterns[3340] = 32'b1001011100110101_1_01_011_101_111_0_x_00;
      patterns[3341] = 32'b1010011100110101_1_10_011_101_111_0_x_00;
      patterns[3342] = 32'b1011011100110101_1_11_011_101_111_0_x_00;
      patterns[3343] = 32'b0101011100110000_1_xx_011_xxx_111_0_1_01;
      patterns[3344] = 32'b0100011100110000_0_xx_011_111_xxx_1_x_xx;
      patterns[3345] = 32'b0000011101101111_1_xx_xxx_xxx_111_0_x_10;
      patterns[3346] = 32'b1000011100110110_1_00_011_110_111_0_x_00;
      patterns[3347] = 32'b1001011100110110_1_01_011_110_111_0_x_00;
      patterns[3348] = 32'b1010011100110110_1_10_011_110_111_0_x_00;
      patterns[3349] = 32'b1011011100110110_1_11_011_110_111_0_x_00;
      patterns[3350] = 32'b0101011100110000_1_xx_011_xxx_111_0_1_01;
      patterns[3351] = 32'b0100011100110000_0_xx_011_111_xxx_1_x_xx;
      patterns[3352] = 32'b0000011100100100_1_xx_xxx_xxx_111_0_x_10;
      patterns[3353] = 32'b1000011100110111_1_00_011_111_111_0_x_00;
      patterns[3354] = 32'b1001011100110111_1_01_011_111_111_0_x_00;
      patterns[3355] = 32'b1010011100110111_1_10_011_111_111_0_x_00;
      patterns[3356] = 32'b1011011100110111_1_11_011_111_111_0_x_00;
      patterns[3357] = 32'b0101011100110000_1_xx_011_xxx_111_0_1_01;
      patterns[3358] = 32'b0100011100110000_0_xx_011_111_xxx_1_x_xx;
      patterns[3359] = 32'b0000011111011100_1_xx_xxx_xxx_111_0_x_10;
      patterns[3360] = 32'b1000011101000000_1_00_100_000_111_0_x_00;
      patterns[3361] = 32'b1001011101000000_1_01_100_000_111_0_x_00;
      patterns[3362] = 32'b1010011101000000_1_10_100_000_111_0_x_00;
      patterns[3363] = 32'b1011011101000000_1_11_100_000_111_0_x_00;
      patterns[3364] = 32'b0101011101000000_1_xx_100_xxx_111_0_1_01;
      patterns[3365] = 32'b0100011101000000_0_xx_100_111_xxx_1_x_xx;
      patterns[3366] = 32'b0000011100001010_1_xx_xxx_xxx_111_0_x_10;
      patterns[3367] = 32'b1000011101000001_1_00_100_001_111_0_x_00;
      patterns[3368] = 32'b1001011101000001_1_01_100_001_111_0_x_00;
      patterns[3369] = 32'b1010011101000001_1_10_100_001_111_0_x_00;
      patterns[3370] = 32'b1011011101000001_1_11_100_001_111_0_x_00;
      patterns[3371] = 32'b0101011101000000_1_xx_100_xxx_111_0_1_01;
      patterns[3372] = 32'b0100011101000000_0_xx_100_111_xxx_1_x_xx;
      patterns[3373] = 32'b0000011100010110_1_xx_xxx_xxx_111_0_x_10;
      patterns[3374] = 32'b1000011101000010_1_00_100_010_111_0_x_00;
      patterns[3375] = 32'b1001011101000010_1_01_100_010_111_0_x_00;
      patterns[3376] = 32'b1010011101000010_1_10_100_010_111_0_x_00;
      patterns[3377] = 32'b1011011101000010_1_11_100_010_111_0_x_00;
      patterns[3378] = 32'b0101011101000000_1_xx_100_xxx_111_0_1_01;
      patterns[3379] = 32'b0100011101000000_0_xx_100_111_xxx_1_x_xx;
      patterns[3380] = 32'b0000011101100011_1_xx_xxx_xxx_111_0_x_10;
      patterns[3381] = 32'b1000011101000011_1_00_100_011_111_0_x_00;
      patterns[3382] = 32'b1001011101000011_1_01_100_011_111_0_x_00;
      patterns[3383] = 32'b1010011101000011_1_10_100_011_111_0_x_00;
      patterns[3384] = 32'b1011011101000011_1_11_100_011_111_0_x_00;
      patterns[3385] = 32'b0101011101000000_1_xx_100_xxx_111_0_1_01;
      patterns[3386] = 32'b0100011101000000_0_xx_100_111_xxx_1_x_xx;
      patterns[3387] = 32'b0000011111101001_1_xx_xxx_xxx_111_0_x_10;
      patterns[3388] = 32'b1000011101000100_1_00_100_100_111_0_x_00;
      patterns[3389] = 32'b1001011101000100_1_01_100_100_111_0_x_00;
      patterns[3390] = 32'b1010011101000100_1_10_100_100_111_0_x_00;
      patterns[3391] = 32'b1011011101000100_1_11_100_100_111_0_x_00;
      patterns[3392] = 32'b0101011101000000_1_xx_100_xxx_111_0_1_01;
      patterns[3393] = 32'b0100011101000000_0_xx_100_111_xxx_1_x_xx;
      patterns[3394] = 32'b0000011110110110_1_xx_xxx_xxx_111_0_x_10;
      patterns[3395] = 32'b1000011101000101_1_00_100_101_111_0_x_00;
      patterns[3396] = 32'b1001011101000101_1_01_100_101_111_0_x_00;
      patterns[3397] = 32'b1010011101000101_1_10_100_101_111_0_x_00;
      patterns[3398] = 32'b1011011101000101_1_11_100_101_111_0_x_00;
      patterns[3399] = 32'b0101011101000000_1_xx_100_xxx_111_0_1_01;
      patterns[3400] = 32'b0100011101000000_0_xx_100_111_xxx_1_x_xx;
      patterns[3401] = 32'b0000011101001001_1_xx_xxx_xxx_111_0_x_10;
      patterns[3402] = 32'b1000011101000110_1_00_100_110_111_0_x_00;
      patterns[3403] = 32'b1001011101000110_1_01_100_110_111_0_x_00;
      patterns[3404] = 32'b1010011101000110_1_10_100_110_111_0_x_00;
      patterns[3405] = 32'b1011011101000110_1_11_100_110_111_0_x_00;
      patterns[3406] = 32'b0101011101000000_1_xx_100_xxx_111_0_1_01;
      patterns[3407] = 32'b0100011101000000_0_xx_100_111_xxx_1_x_xx;
      patterns[3408] = 32'b0000011111101010_1_xx_xxx_xxx_111_0_x_10;
      patterns[3409] = 32'b1000011101000111_1_00_100_111_111_0_x_00;
      patterns[3410] = 32'b1001011101000111_1_01_100_111_111_0_x_00;
      patterns[3411] = 32'b1010011101000111_1_10_100_111_111_0_x_00;
      patterns[3412] = 32'b1011011101000111_1_11_100_111_111_0_x_00;
      patterns[3413] = 32'b0101011101000000_1_xx_100_xxx_111_0_1_01;
      patterns[3414] = 32'b0100011101000000_0_xx_100_111_xxx_1_x_xx;
      patterns[3415] = 32'b0000011100111110_1_xx_xxx_xxx_111_0_x_10;
      patterns[3416] = 32'b1000011101010000_1_00_101_000_111_0_x_00;
      patterns[3417] = 32'b1001011101010000_1_01_101_000_111_0_x_00;
      patterns[3418] = 32'b1010011101010000_1_10_101_000_111_0_x_00;
      patterns[3419] = 32'b1011011101010000_1_11_101_000_111_0_x_00;
      patterns[3420] = 32'b0101011101010000_1_xx_101_xxx_111_0_1_01;
      patterns[3421] = 32'b0100011101010000_0_xx_101_111_xxx_1_x_xx;
      patterns[3422] = 32'b0000011100000110_1_xx_xxx_xxx_111_0_x_10;
      patterns[3423] = 32'b1000011101010001_1_00_101_001_111_0_x_00;
      patterns[3424] = 32'b1001011101010001_1_01_101_001_111_0_x_00;
      patterns[3425] = 32'b1010011101010001_1_10_101_001_111_0_x_00;
      patterns[3426] = 32'b1011011101010001_1_11_101_001_111_0_x_00;
      patterns[3427] = 32'b0101011101010000_1_xx_101_xxx_111_0_1_01;
      patterns[3428] = 32'b0100011101010000_0_xx_101_111_xxx_1_x_xx;
      patterns[3429] = 32'b0000011111001010_1_xx_xxx_xxx_111_0_x_10;
      patterns[3430] = 32'b1000011101010010_1_00_101_010_111_0_x_00;
      patterns[3431] = 32'b1001011101010010_1_01_101_010_111_0_x_00;
      patterns[3432] = 32'b1010011101010010_1_10_101_010_111_0_x_00;
      patterns[3433] = 32'b1011011101010010_1_11_101_010_111_0_x_00;
      patterns[3434] = 32'b0101011101010000_1_xx_101_xxx_111_0_1_01;
      patterns[3435] = 32'b0100011101010000_0_xx_101_111_xxx_1_x_xx;
      patterns[3436] = 32'b0000011100011011_1_xx_xxx_xxx_111_0_x_10;
      patterns[3437] = 32'b1000011101010011_1_00_101_011_111_0_x_00;
      patterns[3438] = 32'b1001011101010011_1_01_101_011_111_0_x_00;
      patterns[3439] = 32'b1010011101010011_1_10_101_011_111_0_x_00;
      patterns[3440] = 32'b1011011101010011_1_11_101_011_111_0_x_00;
      patterns[3441] = 32'b0101011101010000_1_xx_101_xxx_111_0_1_01;
      patterns[3442] = 32'b0100011101010000_0_xx_101_111_xxx_1_x_xx;
      patterns[3443] = 32'b0000011100011010_1_xx_xxx_xxx_111_0_x_10;
      patterns[3444] = 32'b1000011101010100_1_00_101_100_111_0_x_00;
      patterns[3445] = 32'b1001011101010100_1_01_101_100_111_0_x_00;
      patterns[3446] = 32'b1010011101010100_1_10_101_100_111_0_x_00;
      patterns[3447] = 32'b1011011101010100_1_11_101_100_111_0_x_00;
      patterns[3448] = 32'b0101011101010000_1_xx_101_xxx_111_0_1_01;
      patterns[3449] = 32'b0100011101010000_0_xx_101_111_xxx_1_x_xx;
      patterns[3450] = 32'b0000011111000000_1_xx_xxx_xxx_111_0_x_10;
      patterns[3451] = 32'b1000011101010101_1_00_101_101_111_0_x_00;
      patterns[3452] = 32'b1001011101010101_1_01_101_101_111_0_x_00;
      patterns[3453] = 32'b1010011101010101_1_10_101_101_111_0_x_00;
      patterns[3454] = 32'b1011011101010101_1_11_101_101_111_0_x_00;
      patterns[3455] = 32'b0101011101010000_1_xx_101_xxx_111_0_1_01;
      patterns[3456] = 32'b0100011101010000_0_xx_101_111_xxx_1_x_xx;
      patterns[3457] = 32'b0000011100100000_1_xx_xxx_xxx_111_0_x_10;
      patterns[3458] = 32'b1000011101010110_1_00_101_110_111_0_x_00;
      patterns[3459] = 32'b1001011101010110_1_01_101_110_111_0_x_00;
      patterns[3460] = 32'b1010011101010110_1_10_101_110_111_0_x_00;
      patterns[3461] = 32'b1011011101010110_1_11_101_110_111_0_x_00;
      patterns[3462] = 32'b0101011101010000_1_xx_101_xxx_111_0_1_01;
      patterns[3463] = 32'b0100011101010000_0_xx_101_111_xxx_1_x_xx;
      patterns[3464] = 32'b0000011111011011_1_xx_xxx_xxx_111_0_x_10;
      patterns[3465] = 32'b1000011101010111_1_00_101_111_111_0_x_00;
      patterns[3466] = 32'b1001011101010111_1_01_101_111_111_0_x_00;
      patterns[3467] = 32'b1010011101010111_1_10_101_111_111_0_x_00;
      patterns[3468] = 32'b1011011101010111_1_11_101_111_111_0_x_00;
      patterns[3469] = 32'b0101011101010000_1_xx_101_xxx_111_0_1_01;
      patterns[3470] = 32'b0100011101010000_0_xx_101_111_xxx_1_x_xx;
      patterns[3471] = 32'b0000011100000101_1_xx_xxx_xxx_111_0_x_10;
      patterns[3472] = 32'b1000011101100000_1_00_110_000_111_0_x_00;
      patterns[3473] = 32'b1001011101100000_1_01_110_000_111_0_x_00;
      patterns[3474] = 32'b1010011101100000_1_10_110_000_111_0_x_00;
      patterns[3475] = 32'b1011011101100000_1_11_110_000_111_0_x_00;
      patterns[3476] = 32'b0101011101100000_1_xx_110_xxx_111_0_1_01;
      patterns[3477] = 32'b0100011101100000_0_xx_110_111_xxx_1_x_xx;
      patterns[3478] = 32'b0000011101000110_1_xx_xxx_xxx_111_0_x_10;
      patterns[3479] = 32'b1000011101100001_1_00_110_001_111_0_x_00;
      patterns[3480] = 32'b1001011101100001_1_01_110_001_111_0_x_00;
      patterns[3481] = 32'b1010011101100001_1_10_110_001_111_0_x_00;
      patterns[3482] = 32'b1011011101100001_1_11_110_001_111_0_x_00;
      patterns[3483] = 32'b0101011101100000_1_xx_110_xxx_111_0_1_01;
      patterns[3484] = 32'b0100011101100000_0_xx_110_111_xxx_1_x_xx;
      patterns[3485] = 32'b0000011110100010_1_xx_xxx_xxx_111_0_x_10;
      patterns[3486] = 32'b1000011101100010_1_00_110_010_111_0_x_00;
      patterns[3487] = 32'b1001011101100010_1_01_110_010_111_0_x_00;
      patterns[3488] = 32'b1010011101100010_1_10_110_010_111_0_x_00;
      patterns[3489] = 32'b1011011101100010_1_11_110_010_111_0_x_00;
      patterns[3490] = 32'b0101011101100000_1_xx_110_xxx_111_0_1_01;
      patterns[3491] = 32'b0100011101100000_0_xx_110_111_xxx_1_x_xx;
      patterns[3492] = 32'b0000011111010101_1_xx_xxx_xxx_111_0_x_10;
      patterns[3493] = 32'b1000011101100011_1_00_110_011_111_0_x_00;
      patterns[3494] = 32'b1001011101100011_1_01_110_011_111_0_x_00;
      patterns[3495] = 32'b1010011101100011_1_10_110_011_111_0_x_00;
      patterns[3496] = 32'b1011011101100011_1_11_110_011_111_0_x_00;
      patterns[3497] = 32'b0101011101100000_1_xx_110_xxx_111_0_1_01;
      patterns[3498] = 32'b0100011101100000_0_xx_110_111_xxx_1_x_xx;
      patterns[3499] = 32'b0000011110001101_1_xx_xxx_xxx_111_0_x_10;
      patterns[3500] = 32'b1000011101100100_1_00_110_100_111_0_x_00;
      patterns[3501] = 32'b1001011101100100_1_01_110_100_111_0_x_00;
      patterns[3502] = 32'b1010011101100100_1_10_110_100_111_0_x_00;
      patterns[3503] = 32'b1011011101100100_1_11_110_100_111_0_x_00;
      patterns[3504] = 32'b0101011101100000_1_xx_110_xxx_111_0_1_01;
      patterns[3505] = 32'b0100011101100000_0_xx_110_111_xxx_1_x_xx;
      patterns[3506] = 32'b0000011101001001_1_xx_xxx_xxx_111_0_x_10;
      patterns[3507] = 32'b1000011101100101_1_00_110_101_111_0_x_00;
      patterns[3508] = 32'b1001011101100101_1_01_110_101_111_0_x_00;
      patterns[3509] = 32'b1010011101100101_1_10_110_101_111_0_x_00;
      patterns[3510] = 32'b1011011101100101_1_11_110_101_111_0_x_00;
      patterns[3511] = 32'b0101011101100000_1_xx_110_xxx_111_0_1_01;
      patterns[3512] = 32'b0100011101100000_0_xx_110_111_xxx_1_x_xx;
      patterns[3513] = 32'b0000011110001000_1_xx_xxx_xxx_111_0_x_10;
      patterns[3514] = 32'b1000011101100110_1_00_110_110_111_0_x_00;
      patterns[3515] = 32'b1001011101100110_1_01_110_110_111_0_x_00;
      patterns[3516] = 32'b1010011101100110_1_10_110_110_111_0_x_00;
      patterns[3517] = 32'b1011011101100110_1_11_110_110_111_0_x_00;
      patterns[3518] = 32'b0101011101100000_1_xx_110_xxx_111_0_1_01;
      patterns[3519] = 32'b0100011101100000_0_xx_110_111_xxx_1_x_xx;
      patterns[3520] = 32'b0000011100100001_1_xx_xxx_xxx_111_0_x_10;
      patterns[3521] = 32'b1000011101100111_1_00_110_111_111_0_x_00;
      patterns[3522] = 32'b1001011101100111_1_01_110_111_111_0_x_00;
      patterns[3523] = 32'b1010011101100111_1_10_110_111_111_0_x_00;
      patterns[3524] = 32'b1011011101100111_1_11_110_111_111_0_x_00;
      patterns[3525] = 32'b0101011101100000_1_xx_110_xxx_111_0_1_01;
      patterns[3526] = 32'b0100011101100000_0_xx_110_111_xxx_1_x_xx;
      patterns[3527] = 32'b0000011101001011_1_xx_xxx_xxx_111_0_x_10;
      patterns[3528] = 32'b1000011101110000_1_00_111_000_111_0_x_00;
      patterns[3529] = 32'b1001011101110000_1_01_111_000_111_0_x_00;
      patterns[3530] = 32'b1010011101110000_1_10_111_000_111_0_x_00;
      patterns[3531] = 32'b1011011101110000_1_11_111_000_111_0_x_00;
      patterns[3532] = 32'b0101011101110000_1_xx_111_xxx_111_0_1_01;
      patterns[3533] = 32'b0100011101110000_0_xx_111_111_xxx_1_x_xx;
      patterns[3534] = 32'b0000011111011111_1_xx_xxx_xxx_111_0_x_10;
      patterns[3535] = 32'b1000011101110001_1_00_111_001_111_0_x_00;
      patterns[3536] = 32'b1001011101110001_1_01_111_001_111_0_x_00;
      patterns[3537] = 32'b1010011101110001_1_10_111_001_111_0_x_00;
      patterns[3538] = 32'b1011011101110001_1_11_111_001_111_0_x_00;
      patterns[3539] = 32'b0101011101110000_1_xx_111_xxx_111_0_1_01;
      patterns[3540] = 32'b0100011101110000_0_xx_111_111_xxx_1_x_xx;
      patterns[3541] = 32'b0000011110000111_1_xx_xxx_xxx_111_0_x_10;
      patterns[3542] = 32'b1000011101110010_1_00_111_010_111_0_x_00;
      patterns[3543] = 32'b1001011101110010_1_01_111_010_111_0_x_00;
      patterns[3544] = 32'b1010011101110010_1_10_111_010_111_0_x_00;
      patterns[3545] = 32'b1011011101110010_1_11_111_010_111_0_x_00;
      patterns[3546] = 32'b0101011101110000_1_xx_111_xxx_111_0_1_01;
      patterns[3547] = 32'b0100011101110000_0_xx_111_111_xxx_1_x_xx;
      patterns[3548] = 32'b0000011100000110_1_xx_xxx_xxx_111_0_x_10;
      patterns[3549] = 32'b1000011101110011_1_00_111_011_111_0_x_00;
      patterns[3550] = 32'b1001011101110011_1_01_111_011_111_0_x_00;
      patterns[3551] = 32'b1010011101110011_1_10_111_011_111_0_x_00;
      patterns[3552] = 32'b1011011101110011_1_11_111_011_111_0_x_00;
      patterns[3553] = 32'b0101011101110000_1_xx_111_xxx_111_0_1_01;
      patterns[3554] = 32'b0100011101110000_0_xx_111_111_xxx_1_x_xx;
      patterns[3555] = 32'b0000011110000111_1_xx_xxx_xxx_111_0_x_10;
      patterns[3556] = 32'b1000011101110100_1_00_111_100_111_0_x_00;
      patterns[3557] = 32'b1001011101110100_1_01_111_100_111_0_x_00;
      patterns[3558] = 32'b1010011101110100_1_10_111_100_111_0_x_00;
      patterns[3559] = 32'b1011011101110100_1_11_111_100_111_0_x_00;
      patterns[3560] = 32'b0101011101110000_1_xx_111_xxx_111_0_1_01;
      patterns[3561] = 32'b0100011101110000_0_xx_111_111_xxx_1_x_xx;
      patterns[3562] = 32'b0000011110111100_1_xx_xxx_xxx_111_0_x_10;
      patterns[3563] = 32'b1000011101110101_1_00_111_101_111_0_x_00;
      patterns[3564] = 32'b1001011101110101_1_01_111_101_111_0_x_00;
      patterns[3565] = 32'b1010011101110101_1_10_111_101_111_0_x_00;
      patterns[3566] = 32'b1011011101110101_1_11_111_101_111_0_x_00;
      patterns[3567] = 32'b0101011101110000_1_xx_111_xxx_111_0_1_01;
      patterns[3568] = 32'b0100011101110000_0_xx_111_111_xxx_1_x_xx;
      patterns[3569] = 32'b0000011100011001_1_xx_xxx_xxx_111_0_x_10;
      patterns[3570] = 32'b1000011101110110_1_00_111_110_111_0_x_00;
      patterns[3571] = 32'b1001011101110110_1_01_111_110_111_0_x_00;
      patterns[3572] = 32'b1010011101110110_1_10_111_110_111_0_x_00;
      patterns[3573] = 32'b1011011101110110_1_11_111_110_111_0_x_00;
      patterns[3574] = 32'b0101011101110000_1_xx_111_xxx_111_0_1_01;
      patterns[3575] = 32'b0100011101110000_0_xx_111_111_xxx_1_x_xx;
      patterns[3576] = 32'b0000011101111000_1_xx_xxx_xxx_111_0_x_10;
      patterns[3577] = 32'b1000011101110111_1_00_111_111_111_0_x_00;
      patterns[3578] = 32'b1001011101110111_1_01_111_111_111_0_x_00;
      patterns[3579] = 32'b1010011101110111_1_10_111_111_111_0_x_00;
      patterns[3580] = 32'b1011011101110111_1_11_111_111_111_0_x_00;
      patterns[3581] = 32'b0101011101110000_1_xx_111_xxx_111_0_1_01;
      patterns[3582] = 32'b0100011101110000_0_xx_111_111_xxx_1_x_xx;
      patterns[3583] = 32'b0000011101001111_1_xx_xxx_xxx_111_0_x_10;

      for (i = 0; i < 3584; i = i + 1)
      begin
        INST = patterns[i][31:16];
        #10;
        if (patterns[i][15] !== 1'hx)
        begin
          if (WE !== patterns[i][15])
          begin
            $display("%d:WE: (assertion error). Expected %h, found %h", i, patterns[i][15], WE);
            $finish;
          end
        end
        if (patterns[i][14:13] !== 2'hx)
        begin
          if (ALUOP !== patterns[i][14:13])
          begin
            $display("%d:ALUOP: (assertion error). Expected %h, found %h", i, patterns[i][14:13], ALUOP);
            $finish;
          end
        end
        if (patterns[i][12:10] !== 3'hx)
        begin
          if (RS1 !== patterns[i][12:10])
          begin
            $display("%d:RS1: (assertion error). Expected %h, found %h", i, patterns[i][12:10], RS1);
            $finish;
          end
        end
        if (patterns[i][9:7] !== 3'hx)
        begin
          if (RS2 !== patterns[i][9:7])
          begin
            $display("%d:RS2: (assertion error). Expected %h, found %h", i, patterns[i][9:7], RS2);
            $finish;
          end
        end
        if (patterns[i][6:4] !== 3'hx)
        begin
          if (WS !== patterns[i][6:4])
          begin
            $display("%d:WS: (assertion error). Expected %h, found %h", i, patterns[i][6:4], WS);
            $finish;
          end
        end
        if (patterns[i][3] !== 1'hx)
        begin
          if (STR !== patterns[i][3])
          begin
            $display("%d:STR: (assertion error). Expected %h, found %h", i, patterns[i][3], STR);
            $finish;
          end
        end
        if (patterns[i][2] !== 1'hx)
        begin
          if (LDR !== patterns[i][2])
          begin
            $display("%d:LDR: (assertion error). Expected %h, found %h", i, patterns[i][2], LDR);
            $finish;
          end
        end
        if (patterns[i][1:0] !== 2'hx)
        begin
          if (DMUX !== patterns[i][1:0])
          begin
            $display("%d:DMUX: (assertion error). Expected %h, found %h", i, patterns[i][1:0], DMUX);
            $finish;
          end
        end
      end

      $display("All tests passed.");
    end
    endmodule
