--  A testbench for control_unit_ALUOP_tb
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity control_unit_ALUOP_tb is
end control_unit_ALUOP_tb;

architecture behav of control_unit_ALUOP_tb is
  component main
    port (
      INST: in std_logic_vector(15 downto 0);
      FL_Z: in std_logic;
      ALUOP: out std_logic_vector(1 downto 0);
      RS1: out std_logic_vector(2 downto 0);
      RS2: out std_logic_vector(2 downto 0);
      WS: out std_logic_vector(2 downto 0);
      STR: out std_logic;
      WE: out std_logic;
      DMUX: out std_logic_vector(1 downto 0);
      LDR: out std_logic;
      FL_EN: out std_logic;
      HE: out std_logic);
  end component;

  signal INST : std_logic_vector(15 downto 0);
  signal FL_Z : std_logic;
  signal ALUOP : std_logic_vector(1 downto 0);
  signal RS1 : std_logic_vector(2 downto 0);
  signal RS2 : std_logic_vector(2 downto 0);
  signal WS : std_logic_vector(2 downto 0);
  signal STR : std_logic;
  signal WE : std_logic;
  signal DMUX : std_logic_vector(1 downto 0);
  signal LDR : std_logic;
  signal FL_EN : std_logic;
  signal HE : std_logic;
  function to_string ( a: std_logic_vector) return string is
      variable b : string (1 to a'length) := (others => NUL);
      variable stri : integer := 1; 
  begin
      for i in a'range loop
          b(stri) := std_logic'image(a((i)))(2);
      stri := stri+1;
      end loop;
      return b;
  end function;
begin
  main_0 : main port map (
    INST => INST,
    FL_Z => FL_Z,
    ALUOP => ALUOP,
    RS1 => RS1,
    RS2 => RS2,
    WS => WS,
    STR => STR,
    WE => WE,
    DMUX => DMUX,
    LDR => LDR,
    FL_EN => FL_EN,
    HE => HE );
  process
    type pattern_type is record
      INST : std_logic_vector(15 downto 0);
      ALUOP : std_logic_vector(1 downto 0);
    end record;
    type pattern_array is array (natural range <>) of pattern_type;
    constant patterns : pattern_array := (
      ("1000000000000000", "00"), -- i=0
      ("1001000000000000", "01"), -- i=1
      ("1010000000000000", "10"), -- i=2
      ("1011000000000000", "11"), -- i=3
      ("1000000000000001", "00"), -- i=4
      ("1001000000000001", "01"), -- i=5
      ("1010000000000001", "10"), -- i=6
      ("1011000000000001", "11"), -- i=7
      ("1000000000000010", "00"), -- i=8
      ("1001000000000010", "01"), -- i=9
      ("1010000000000010", "10"), -- i=10
      ("1011000000000010", "11"), -- i=11
      ("1000000000000011", "00"), -- i=12
      ("1001000000000011", "01"), -- i=13
      ("1010000000000011", "10"), -- i=14
      ("1011000000000011", "11"), -- i=15
      ("1000000000000100", "00"), -- i=16
      ("1001000000000100", "01"), -- i=17
      ("1010000000000100", "10"), -- i=18
      ("1011000000000100", "11"), -- i=19
      ("1000000000000101", "00"), -- i=20
      ("1001000000000101", "01"), -- i=21
      ("1010000000000101", "10"), -- i=22
      ("1011000000000101", "11"), -- i=23
      ("1000000000000110", "00"), -- i=24
      ("1001000000000110", "01"), -- i=25
      ("1010000000000110", "10"), -- i=26
      ("1011000000000110", "11"), -- i=27
      ("1000000000000111", "00"), -- i=28
      ("1001000000000111", "01"), -- i=29
      ("1010000000000111", "10"), -- i=30
      ("1011000000000111", "11"), -- i=31
      ("1000000000010000", "00"), -- i=32
      ("1001000000010000", "01"), -- i=33
      ("1010000000010000", "10"), -- i=34
      ("1011000000010000", "11"), -- i=35
      ("1000000000010001", "00"), -- i=36
      ("1001000000010001", "01"), -- i=37
      ("1010000000010001", "10"), -- i=38
      ("1011000000010001", "11"), -- i=39
      ("1000000000010010", "00"), -- i=40
      ("1001000000010010", "01"), -- i=41
      ("1010000000010010", "10"), -- i=42
      ("1011000000010010", "11"), -- i=43
      ("1000000000010011", "00"), -- i=44
      ("1001000000010011", "01"), -- i=45
      ("1010000000010011", "10"), -- i=46
      ("1011000000010011", "11"), -- i=47
      ("1000000000010100", "00"), -- i=48
      ("1001000000010100", "01"), -- i=49
      ("1010000000010100", "10"), -- i=50
      ("1011000000010100", "11"), -- i=51
      ("1000000000010101", "00"), -- i=52
      ("1001000000010101", "01"), -- i=53
      ("1010000000010101", "10"), -- i=54
      ("1011000000010101", "11"), -- i=55
      ("1000000000010110", "00"), -- i=56
      ("1001000000010110", "01"), -- i=57
      ("1010000000010110", "10"), -- i=58
      ("1011000000010110", "11"), -- i=59
      ("1000000000010111", "00"), -- i=60
      ("1001000000010111", "01"), -- i=61
      ("1010000000010111", "10"), -- i=62
      ("1011000000010111", "11"), -- i=63
      ("1000000000100000", "00"), -- i=64
      ("1001000000100000", "01"), -- i=65
      ("1010000000100000", "10"), -- i=66
      ("1011000000100000", "11"), -- i=67
      ("1000000000100001", "00"), -- i=68
      ("1001000000100001", "01"), -- i=69
      ("1010000000100001", "10"), -- i=70
      ("1011000000100001", "11"), -- i=71
      ("1000000000100010", "00"), -- i=72
      ("1001000000100010", "01"), -- i=73
      ("1010000000100010", "10"), -- i=74
      ("1011000000100010", "11"), -- i=75
      ("1000000000100011", "00"), -- i=76
      ("1001000000100011", "01"), -- i=77
      ("1010000000100011", "10"), -- i=78
      ("1011000000100011", "11"), -- i=79
      ("1000000000100100", "00"), -- i=80
      ("1001000000100100", "01"), -- i=81
      ("1010000000100100", "10"), -- i=82
      ("1011000000100100", "11"), -- i=83
      ("1000000000100101", "00"), -- i=84
      ("1001000000100101", "01"), -- i=85
      ("1010000000100101", "10"), -- i=86
      ("1011000000100101", "11"), -- i=87
      ("1000000000100110", "00"), -- i=88
      ("1001000000100110", "01"), -- i=89
      ("1010000000100110", "10"), -- i=90
      ("1011000000100110", "11"), -- i=91
      ("1000000000100111", "00"), -- i=92
      ("1001000000100111", "01"), -- i=93
      ("1010000000100111", "10"), -- i=94
      ("1011000000100111", "11"), -- i=95
      ("1000000000110000", "00"), -- i=96
      ("1001000000110000", "01"), -- i=97
      ("1010000000110000", "10"), -- i=98
      ("1011000000110000", "11"), -- i=99
      ("1000000000110001", "00"), -- i=100
      ("1001000000110001", "01"), -- i=101
      ("1010000000110001", "10"), -- i=102
      ("1011000000110001", "11"), -- i=103
      ("1000000000110010", "00"), -- i=104
      ("1001000000110010", "01"), -- i=105
      ("1010000000110010", "10"), -- i=106
      ("1011000000110010", "11"), -- i=107
      ("1000000000110011", "00"), -- i=108
      ("1001000000110011", "01"), -- i=109
      ("1010000000110011", "10"), -- i=110
      ("1011000000110011", "11"), -- i=111
      ("1000000000110100", "00"), -- i=112
      ("1001000000110100", "01"), -- i=113
      ("1010000000110100", "10"), -- i=114
      ("1011000000110100", "11"), -- i=115
      ("1000000000110101", "00"), -- i=116
      ("1001000000110101", "01"), -- i=117
      ("1010000000110101", "10"), -- i=118
      ("1011000000110101", "11"), -- i=119
      ("1000000000110110", "00"), -- i=120
      ("1001000000110110", "01"), -- i=121
      ("1010000000110110", "10"), -- i=122
      ("1011000000110110", "11"), -- i=123
      ("1000000000110111", "00"), -- i=124
      ("1001000000110111", "01"), -- i=125
      ("1010000000110111", "10"), -- i=126
      ("1011000000110111", "11"), -- i=127
      ("1000000001000000", "00"), -- i=128
      ("1001000001000000", "01"), -- i=129
      ("1010000001000000", "10"), -- i=130
      ("1011000001000000", "11"), -- i=131
      ("1000000001000001", "00"), -- i=132
      ("1001000001000001", "01"), -- i=133
      ("1010000001000001", "10"), -- i=134
      ("1011000001000001", "11"), -- i=135
      ("1000000001000010", "00"), -- i=136
      ("1001000001000010", "01"), -- i=137
      ("1010000001000010", "10"), -- i=138
      ("1011000001000010", "11"), -- i=139
      ("1000000001000011", "00"), -- i=140
      ("1001000001000011", "01"), -- i=141
      ("1010000001000011", "10"), -- i=142
      ("1011000001000011", "11"), -- i=143
      ("1000000001000100", "00"), -- i=144
      ("1001000001000100", "01"), -- i=145
      ("1010000001000100", "10"), -- i=146
      ("1011000001000100", "11"), -- i=147
      ("1000000001000101", "00"), -- i=148
      ("1001000001000101", "01"), -- i=149
      ("1010000001000101", "10"), -- i=150
      ("1011000001000101", "11"), -- i=151
      ("1000000001000110", "00"), -- i=152
      ("1001000001000110", "01"), -- i=153
      ("1010000001000110", "10"), -- i=154
      ("1011000001000110", "11"), -- i=155
      ("1000000001000111", "00"), -- i=156
      ("1001000001000111", "01"), -- i=157
      ("1010000001000111", "10"), -- i=158
      ("1011000001000111", "11"), -- i=159
      ("1000000001010000", "00"), -- i=160
      ("1001000001010000", "01"), -- i=161
      ("1010000001010000", "10"), -- i=162
      ("1011000001010000", "11"), -- i=163
      ("1000000001010001", "00"), -- i=164
      ("1001000001010001", "01"), -- i=165
      ("1010000001010001", "10"), -- i=166
      ("1011000001010001", "11"), -- i=167
      ("1000000001010010", "00"), -- i=168
      ("1001000001010010", "01"), -- i=169
      ("1010000001010010", "10"), -- i=170
      ("1011000001010010", "11"), -- i=171
      ("1000000001010011", "00"), -- i=172
      ("1001000001010011", "01"), -- i=173
      ("1010000001010011", "10"), -- i=174
      ("1011000001010011", "11"), -- i=175
      ("1000000001010100", "00"), -- i=176
      ("1001000001010100", "01"), -- i=177
      ("1010000001010100", "10"), -- i=178
      ("1011000001010100", "11"), -- i=179
      ("1000000001010101", "00"), -- i=180
      ("1001000001010101", "01"), -- i=181
      ("1010000001010101", "10"), -- i=182
      ("1011000001010101", "11"), -- i=183
      ("1000000001010110", "00"), -- i=184
      ("1001000001010110", "01"), -- i=185
      ("1010000001010110", "10"), -- i=186
      ("1011000001010110", "11"), -- i=187
      ("1000000001010111", "00"), -- i=188
      ("1001000001010111", "01"), -- i=189
      ("1010000001010111", "10"), -- i=190
      ("1011000001010111", "11"), -- i=191
      ("1000000001100000", "00"), -- i=192
      ("1001000001100000", "01"), -- i=193
      ("1010000001100000", "10"), -- i=194
      ("1011000001100000", "11"), -- i=195
      ("1000000001100001", "00"), -- i=196
      ("1001000001100001", "01"), -- i=197
      ("1010000001100001", "10"), -- i=198
      ("1011000001100001", "11"), -- i=199
      ("1000000001100010", "00"), -- i=200
      ("1001000001100010", "01"), -- i=201
      ("1010000001100010", "10"), -- i=202
      ("1011000001100010", "11"), -- i=203
      ("1000000001100011", "00"), -- i=204
      ("1001000001100011", "01"), -- i=205
      ("1010000001100011", "10"), -- i=206
      ("1011000001100011", "11"), -- i=207
      ("1000000001100100", "00"), -- i=208
      ("1001000001100100", "01"), -- i=209
      ("1010000001100100", "10"), -- i=210
      ("1011000001100100", "11"), -- i=211
      ("1000000001100101", "00"), -- i=212
      ("1001000001100101", "01"), -- i=213
      ("1010000001100101", "10"), -- i=214
      ("1011000001100101", "11"), -- i=215
      ("1000000001100110", "00"), -- i=216
      ("1001000001100110", "01"), -- i=217
      ("1010000001100110", "10"), -- i=218
      ("1011000001100110", "11"), -- i=219
      ("1000000001100111", "00"), -- i=220
      ("1001000001100111", "01"), -- i=221
      ("1010000001100111", "10"), -- i=222
      ("1011000001100111", "11"), -- i=223
      ("1000000001110000", "00"), -- i=224
      ("1001000001110000", "01"), -- i=225
      ("1010000001110000", "10"), -- i=226
      ("1011000001110000", "11"), -- i=227
      ("1000000001110001", "00"), -- i=228
      ("1001000001110001", "01"), -- i=229
      ("1010000001110001", "10"), -- i=230
      ("1011000001110001", "11"), -- i=231
      ("1000000001110010", "00"), -- i=232
      ("1001000001110010", "01"), -- i=233
      ("1010000001110010", "10"), -- i=234
      ("1011000001110010", "11"), -- i=235
      ("1000000001110011", "00"), -- i=236
      ("1001000001110011", "01"), -- i=237
      ("1010000001110011", "10"), -- i=238
      ("1011000001110011", "11"), -- i=239
      ("1000000001110100", "00"), -- i=240
      ("1001000001110100", "01"), -- i=241
      ("1010000001110100", "10"), -- i=242
      ("1011000001110100", "11"), -- i=243
      ("1000000001110101", "00"), -- i=244
      ("1001000001110101", "01"), -- i=245
      ("1010000001110101", "10"), -- i=246
      ("1011000001110101", "11"), -- i=247
      ("1000000001110110", "00"), -- i=248
      ("1001000001110110", "01"), -- i=249
      ("1010000001110110", "10"), -- i=250
      ("1011000001110110", "11"), -- i=251
      ("1000000001110111", "00"), -- i=252
      ("1001000001110111", "01"), -- i=253
      ("1010000001110111", "10"), -- i=254
      ("1011000001110111", "11"), -- i=255
      ("1000000100000000", "00"), -- i=256
      ("1001000100000000", "01"), -- i=257
      ("1010000100000000", "10"), -- i=258
      ("1011000100000000", "11"), -- i=259
      ("1000000100000001", "00"), -- i=260
      ("1001000100000001", "01"), -- i=261
      ("1010000100000001", "10"), -- i=262
      ("1011000100000001", "11"), -- i=263
      ("1000000100000010", "00"), -- i=264
      ("1001000100000010", "01"), -- i=265
      ("1010000100000010", "10"), -- i=266
      ("1011000100000010", "11"), -- i=267
      ("1000000100000011", "00"), -- i=268
      ("1001000100000011", "01"), -- i=269
      ("1010000100000011", "10"), -- i=270
      ("1011000100000011", "11"), -- i=271
      ("1000000100000100", "00"), -- i=272
      ("1001000100000100", "01"), -- i=273
      ("1010000100000100", "10"), -- i=274
      ("1011000100000100", "11"), -- i=275
      ("1000000100000101", "00"), -- i=276
      ("1001000100000101", "01"), -- i=277
      ("1010000100000101", "10"), -- i=278
      ("1011000100000101", "11"), -- i=279
      ("1000000100000110", "00"), -- i=280
      ("1001000100000110", "01"), -- i=281
      ("1010000100000110", "10"), -- i=282
      ("1011000100000110", "11"), -- i=283
      ("1000000100000111", "00"), -- i=284
      ("1001000100000111", "01"), -- i=285
      ("1010000100000111", "10"), -- i=286
      ("1011000100000111", "11"), -- i=287
      ("1000000100010000", "00"), -- i=288
      ("1001000100010000", "01"), -- i=289
      ("1010000100010000", "10"), -- i=290
      ("1011000100010000", "11"), -- i=291
      ("1000000100010001", "00"), -- i=292
      ("1001000100010001", "01"), -- i=293
      ("1010000100010001", "10"), -- i=294
      ("1011000100010001", "11"), -- i=295
      ("1000000100010010", "00"), -- i=296
      ("1001000100010010", "01"), -- i=297
      ("1010000100010010", "10"), -- i=298
      ("1011000100010010", "11"), -- i=299
      ("1000000100010011", "00"), -- i=300
      ("1001000100010011", "01"), -- i=301
      ("1010000100010011", "10"), -- i=302
      ("1011000100010011", "11"), -- i=303
      ("1000000100010100", "00"), -- i=304
      ("1001000100010100", "01"), -- i=305
      ("1010000100010100", "10"), -- i=306
      ("1011000100010100", "11"), -- i=307
      ("1000000100010101", "00"), -- i=308
      ("1001000100010101", "01"), -- i=309
      ("1010000100010101", "10"), -- i=310
      ("1011000100010101", "11"), -- i=311
      ("1000000100010110", "00"), -- i=312
      ("1001000100010110", "01"), -- i=313
      ("1010000100010110", "10"), -- i=314
      ("1011000100010110", "11"), -- i=315
      ("1000000100010111", "00"), -- i=316
      ("1001000100010111", "01"), -- i=317
      ("1010000100010111", "10"), -- i=318
      ("1011000100010111", "11"), -- i=319
      ("1000000100100000", "00"), -- i=320
      ("1001000100100000", "01"), -- i=321
      ("1010000100100000", "10"), -- i=322
      ("1011000100100000", "11"), -- i=323
      ("1000000100100001", "00"), -- i=324
      ("1001000100100001", "01"), -- i=325
      ("1010000100100001", "10"), -- i=326
      ("1011000100100001", "11"), -- i=327
      ("1000000100100010", "00"), -- i=328
      ("1001000100100010", "01"), -- i=329
      ("1010000100100010", "10"), -- i=330
      ("1011000100100010", "11"), -- i=331
      ("1000000100100011", "00"), -- i=332
      ("1001000100100011", "01"), -- i=333
      ("1010000100100011", "10"), -- i=334
      ("1011000100100011", "11"), -- i=335
      ("1000000100100100", "00"), -- i=336
      ("1001000100100100", "01"), -- i=337
      ("1010000100100100", "10"), -- i=338
      ("1011000100100100", "11"), -- i=339
      ("1000000100100101", "00"), -- i=340
      ("1001000100100101", "01"), -- i=341
      ("1010000100100101", "10"), -- i=342
      ("1011000100100101", "11"), -- i=343
      ("1000000100100110", "00"), -- i=344
      ("1001000100100110", "01"), -- i=345
      ("1010000100100110", "10"), -- i=346
      ("1011000100100110", "11"), -- i=347
      ("1000000100100111", "00"), -- i=348
      ("1001000100100111", "01"), -- i=349
      ("1010000100100111", "10"), -- i=350
      ("1011000100100111", "11"), -- i=351
      ("1000000100110000", "00"), -- i=352
      ("1001000100110000", "01"), -- i=353
      ("1010000100110000", "10"), -- i=354
      ("1011000100110000", "11"), -- i=355
      ("1000000100110001", "00"), -- i=356
      ("1001000100110001", "01"), -- i=357
      ("1010000100110001", "10"), -- i=358
      ("1011000100110001", "11"), -- i=359
      ("1000000100110010", "00"), -- i=360
      ("1001000100110010", "01"), -- i=361
      ("1010000100110010", "10"), -- i=362
      ("1011000100110010", "11"), -- i=363
      ("1000000100110011", "00"), -- i=364
      ("1001000100110011", "01"), -- i=365
      ("1010000100110011", "10"), -- i=366
      ("1011000100110011", "11"), -- i=367
      ("1000000100110100", "00"), -- i=368
      ("1001000100110100", "01"), -- i=369
      ("1010000100110100", "10"), -- i=370
      ("1011000100110100", "11"), -- i=371
      ("1000000100110101", "00"), -- i=372
      ("1001000100110101", "01"), -- i=373
      ("1010000100110101", "10"), -- i=374
      ("1011000100110101", "11"), -- i=375
      ("1000000100110110", "00"), -- i=376
      ("1001000100110110", "01"), -- i=377
      ("1010000100110110", "10"), -- i=378
      ("1011000100110110", "11"), -- i=379
      ("1000000100110111", "00"), -- i=380
      ("1001000100110111", "01"), -- i=381
      ("1010000100110111", "10"), -- i=382
      ("1011000100110111", "11"), -- i=383
      ("1000000101000000", "00"), -- i=384
      ("1001000101000000", "01"), -- i=385
      ("1010000101000000", "10"), -- i=386
      ("1011000101000000", "11"), -- i=387
      ("1000000101000001", "00"), -- i=388
      ("1001000101000001", "01"), -- i=389
      ("1010000101000001", "10"), -- i=390
      ("1011000101000001", "11"), -- i=391
      ("1000000101000010", "00"), -- i=392
      ("1001000101000010", "01"), -- i=393
      ("1010000101000010", "10"), -- i=394
      ("1011000101000010", "11"), -- i=395
      ("1000000101000011", "00"), -- i=396
      ("1001000101000011", "01"), -- i=397
      ("1010000101000011", "10"), -- i=398
      ("1011000101000011", "11"), -- i=399
      ("1000000101000100", "00"), -- i=400
      ("1001000101000100", "01"), -- i=401
      ("1010000101000100", "10"), -- i=402
      ("1011000101000100", "11"), -- i=403
      ("1000000101000101", "00"), -- i=404
      ("1001000101000101", "01"), -- i=405
      ("1010000101000101", "10"), -- i=406
      ("1011000101000101", "11"), -- i=407
      ("1000000101000110", "00"), -- i=408
      ("1001000101000110", "01"), -- i=409
      ("1010000101000110", "10"), -- i=410
      ("1011000101000110", "11"), -- i=411
      ("1000000101000111", "00"), -- i=412
      ("1001000101000111", "01"), -- i=413
      ("1010000101000111", "10"), -- i=414
      ("1011000101000111", "11"), -- i=415
      ("1000000101010000", "00"), -- i=416
      ("1001000101010000", "01"), -- i=417
      ("1010000101010000", "10"), -- i=418
      ("1011000101010000", "11"), -- i=419
      ("1000000101010001", "00"), -- i=420
      ("1001000101010001", "01"), -- i=421
      ("1010000101010001", "10"), -- i=422
      ("1011000101010001", "11"), -- i=423
      ("1000000101010010", "00"), -- i=424
      ("1001000101010010", "01"), -- i=425
      ("1010000101010010", "10"), -- i=426
      ("1011000101010010", "11"), -- i=427
      ("1000000101010011", "00"), -- i=428
      ("1001000101010011", "01"), -- i=429
      ("1010000101010011", "10"), -- i=430
      ("1011000101010011", "11"), -- i=431
      ("1000000101010100", "00"), -- i=432
      ("1001000101010100", "01"), -- i=433
      ("1010000101010100", "10"), -- i=434
      ("1011000101010100", "11"), -- i=435
      ("1000000101010101", "00"), -- i=436
      ("1001000101010101", "01"), -- i=437
      ("1010000101010101", "10"), -- i=438
      ("1011000101010101", "11"), -- i=439
      ("1000000101010110", "00"), -- i=440
      ("1001000101010110", "01"), -- i=441
      ("1010000101010110", "10"), -- i=442
      ("1011000101010110", "11"), -- i=443
      ("1000000101010111", "00"), -- i=444
      ("1001000101010111", "01"), -- i=445
      ("1010000101010111", "10"), -- i=446
      ("1011000101010111", "11"), -- i=447
      ("1000000101100000", "00"), -- i=448
      ("1001000101100000", "01"), -- i=449
      ("1010000101100000", "10"), -- i=450
      ("1011000101100000", "11"), -- i=451
      ("1000000101100001", "00"), -- i=452
      ("1001000101100001", "01"), -- i=453
      ("1010000101100001", "10"), -- i=454
      ("1011000101100001", "11"), -- i=455
      ("1000000101100010", "00"), -- i=456
      ("1001000101100010", "01"), -- i=457
      ("1010000101100010", "10"), -- i=458
      ("1011000101100010", "11"), -- i=459
      ("1000000101100011", "00"), -- i=460
      ("1001000101100011", "01"), -- i=461
      ("1010000101100011", "10"), -- i=462
      ("1011000101100011", "11"), -- i=463
      ("1000000101100100", "00"), -- i=464
      ("1001000101100100", "01"), -- i=465
      ("1010000101100100", "10"), -- i=466
      ("1011000101100100", "11"), -- i=467
      ("1000000101100101", "00"), -- i=468
      ("1001000101100101", "01"), -- i=469
      ("1010000101100101", "10"), -- i=470
      ("1011000101100101", "11"), -- i=471
      ("1000000101100110", "00"), -- i=472
      ("1001000101100110", "01"), -- i=473
      ("1010000101100110", "10"), -- i=474
      ("1011000101100110", "11"), -- i=475
      ("1000000101100111", "00"), -- i=476
      ("1001000101100111", "01"), -- i=477
      ("1010000101100111", "10"), -- i=478
      ("1011000101100111", "11"), -- i=479
      ("1000000101110000", "00"), -- i=480
      ("1001000101110000", "01"), -- i=481
      ("1010000101110000", "10"), -- i=482
      ("1011000101110000", "11"), -- i=483
      ("1000000101110001", "00"), -- i=484
      ("1001000101110001", "01"), -- i=485
      ("1010000101110001", "10"), -- i=486
      ("1011000101110001", "11"), -- i=487
      ("1000000101110010", "00"), -- i=488
      ("1001000101110010", "01"), -- i=489
      ("1010000101110010", "10"), -- i=490
      ("1011000101110010", "11"), -- i=491
      ("1000000101110011", "00"), -- i=492
      ("1001000101110011", "01"), -- i=493
      ("1010000101110011", "10"), -- i=494
      ("1011000101110011", "11"), -- i=495
      ("1000000101110100", "00"), -- i=496
      ("1001000101110100", "01"), -- i=497
      ("1010000101110100", "10"), -- i=498
      ("1011000101110100", "11"), -- i=499
      ("1000000101110101", "00"), -- i=500
      ("1001000101110101", "01"), -- i=501
      ("1010000101110101", "10"), -- i=502
      ("1011000101110101", "11"), -- i=503
      ("1000000101110110", "00"), -- i=504
      ("1001000101110110", "01"), -- i=505
      ("1010000101110110", "10"), -- i=506
      ("1011000101110110", "11"), -- i=507
      ("1000000101110111", "00"), -- i=508
      ("1001000101110111", "01"), -- i=509
      ("1010000101110111", "10"), -- i=510
      ("1011000101110111", "11"), -- i=511
      ("1000001000000000", "00"), -- i=512
      ("1001001000000000", "01"), -- i=513
      ("1010001000000000", "10"), -- i=514
      ("1011001000000000", "11"), -- i=515
      ("1000001000000001", "00"), -- i=516
      ("1001001000000001", "01"), -- i=517
      ("1010001000000001", "10"), -- i=518
      ("1011001000000001", "11"), -- i=519
      ("1000001000000010", "00"), -- i=520
      ("1001001000000010", "01"), -- i=521
      ("1010001000000010", "10"), -- i=522
      ("1011001000000010", "11"), -- i=523
      ("1000001000000011", "00"), -- i=524
      ("1001001000000011", "01"), -- i=525
      ("1010001000000011", "10"), -- i=526
      ("1011001000000011", "11"), -- i=527
      ("1000001000000100", "00"), -- i=528
      ("1001001000000100", "01"), -- i=529
      ("1010001000000100", "10"), -- i=530
      ("1011001000000100", "11"), -- i=531
      ("1000001000000101", "00"), -- i=532
      ("1001001000000101", "01"), -- i=533
      ("1010001000000101", "10"), -- i=534
      ("1011001000000101", "11"), -- i=535
      ("1000001000000110", "00"), -- i=536
      ("1001001000000110", "01"), -- i=537
      ("1010001000000110", "10"), -- i=538
      ("1011001000000110", "11"), -- i=539
      ("1000001000000111", "00"), -- i=540
      ("1001001000000111", "01"), -- i=541
      ("1010001000000111", "10"), -- i=542
      ("1011001000000111", "11"), -- i=543
      ("1000001000010000", "00"), -- i=544
      ("1001001000010000", "01"), -- i=545
      ("1010001000010000", "10"), -- i=546
      ("1011001000010000", "11"), -- i=547
      ("1000001000010001", "00"), -- i=548
      ("1001001000010001", "01"), -- i=549
      ("1010001000010001", "10"), -- i=550
      ("1011001000010001", "11"), -- i=551
      ("1000001000010010", "00"), -- i=552
      ("1001001000010010", "01"), -- i=553
      ("1010001000010010", "10"), -- i=554
      ("1011001000010010", "11"), -- i=555
      ("1000001000010011", "00"), -- i=556
      ("1001001000010011", "01"), -- i=557
      ("1010001000010011", "10"), -- i=558
      ("1011001000010011", "11"), -- i=559
      ("1000001000010100", "00"), -- i=560
      ("1001001000010100", "01"), -- i=561
      ("1010001000010100", "10"), -- i=562
      ("1011001000010100", "11"), -- i=563
      ("1000001000010101", "00"), -- i=564
      ("1001001000010101", "01"), -- i=565
      ("1010001000010101", "10"), -- i=566
      ("1011001000010101", "11"), -- i=567
      ("1000001000010110", "00"), -- i=568
      ("1001001000010110", "01"), -- i=569
      ("1010001000010110", "10"), -- i=570
      ("1011001000010110", "11"), -- i=571
      ("1000001000010111", "00"), -- i=572
      ("1001001000010111", "01"), -- i=573
      ("1010001000010111", "10"), -- i=574
      ("1011001000010111", "11"), -- i=575
      ("1000001000100000", "00"), -- i=576
      ("1001001000100000", "01"), -- i=577
      ("1010001000100000", "10"), -- i=578
      ("1011001000100000", "11"), -- i=579
      ("1000001000100001", "00"), -- i=580
      ("1001001000100001", "01"), -- i=581
      ("1010001000100001", "10"), -- i=582
      ("1011001000100001", "11"), -- i=583
      ("1000001000100010", "00"), -- i=584
      ("1001001000100010", "01"), -- i=585
      ("1010001000100010", "10"), -- i=586
      ("1011001000100010", "11"), -- i=587
      ("1000001000100011", "00"), -- i=588
      ("1001001000100011", "01"), -- i=589
      ("1010001000100011", "10"), -- i=590
      ("1011001000100011", "11"), -- i=591
      ("1000001000100100", "00"), -- i=592
      ("1001001000100100", "01"), -- i=593
      ("1010001000100100", "10"), -- i=594
      ("1011001000100100", "11"), -- i=595
      ("1000001000100101", "00"), -- i=596
      ("1001001000100101", "01"), -- i=597
      ("1010001000100101", "10"), -- i=598
      ("1011001000100101", "11"), -- i=599
      ("1000001000100110", "00"), -- i=600
      ("1001001000100110", "01"), -- i=601
      ("1010001000100110", "10"), -- i=602
      ("1011001000100110", "11"), -- i=603
      ("1000001000100111", "00"), -- i=604
      ("1001001000100111", "01"), -- i=605
      ("1010001000100111", "10"), -- i=606
      ("1011001000100111", "11"), -- i=607
      ("1000001000110000", "00"), -- i=608
      ("1001001000110000", "01"), -- i=609
      ("1010001000110000", "10"), -- i=610
      ("1011001000110000", "11"), -- i=611
      ("1000001000110001", "00"), -- i=612
      ("1001001000110001", "01"), -- i=613
      ("1010001000110001", "10"), -- i=614
      ("1011001000110001", "11"), -- i=615
      ("1000001000110010", "00"), -- i=616
      ("1001001000110010", "01"), -- i=617
      ("1010001000110010", "10"), -- i=618
      ("1011001000110010", "11"), -- i=619
      ("1000001000110011", "00"), -- i=620
      ("1001001000110011", "01"), -- i=621
      ("1010001000110011", "10"), -- i=622
      ("1011001000110011", "11"), -- i=623
      ("1000001000110100", "00"), -- i=624
      ("1001001000110100", "01"), -- i=625
      ("1010001000110100", "10"), -- i=626
      ("1011001000110100", "11"), -- i=627
      ("1000001000110101", "00"), -- i=628
      ("1001001000110101", "01"), -- i=629
      ("1010001000110101", "10"), -- i=630
      ("1011001000110101", "11"), -- i=631
      ("1000001000110110", "00"), -- i=632
      ("1001001000110110", "01"), -- i=633
      ("1010001000110110", "10"), -- i=634
      ("1011001000110110", "11"), -- i=635
      ("1000001000110111", "00"), -- i=636
      ("1001001000110111", "01"), -- i=637
      ("1010001000110111", "10"), -- i=638
      ("1011001000110111", "11"), -- i=639
      ("1000001001000000", "00"), -- i=640
      ("1001001001000000", "01"), -- i=641
      ("1010001001000000", "10"), -- i=642
      ("1011001001000000", "11"), -- i=643
      ("1000001001000001", "00"), -- i=644
      ("1001001001000001", "01"), -- i=645
      ("1010001001000001", "10"), -- i=646
      ("1011001001000001", "11"), -- i=647
      ("1000001001000010", "00"), -- i=648
      ("1001001001000010", "01"), -- i=649
      ("1010001001000010", "10"), -- i=650
      ("1011001001000010", "11"), -- i=651
      ("1000001001000011", "00"), -- i=652
      ("1001001001000011", "01"), -- i=653
      ("1010001001000011", "10"), -- i=654
      ("1011001001000011", "11"), -- i=655
      ("1000001001000100", "00"), -- i=656
      ("1001001001000100", "01"), -- i=657
      ("1010001001000100", "10"), -- i=658
      ("1011001001000100", "11"), -- i=659
      ("1000001001000101", "00"), -- i=660
      ("1001001001000101", "01"), -- i=661
      ("1010001001000101", "10"), -- i=662
      ("1011001001000101", "11"), -- i=663
      ("1000001001000110", "00"), -- i=664
      ("1001001001000110", "01"), -- i=665
      ("1010001001000110", "10"), -- i=666
      ("1011001001000110", "11"), -- i=667
      ("1000001001000111", "00"), -- i=668
      ("1001001001000111", "01"), -- i=669
      ("1010001001000111", "10"), -- i=670
      ("1011001001000111", "11"), -- i=671
      ("1000001001010000", "00"), -- i=672
      ("1001001001010000", "01"), -- i=673
      ("1010001001010000", "10"), -- i=674
      ("1011001001010000", "11"), -- i=675
      ("1000001001010001", "00"), -- i=676
      ("1001001001010001", "01"), -- i=677
      ("1010001001010001", "10"), -- i=678
      ("1011001001010001", "11"), -- i=679
      ("1000001001010010", "00"), -- i=680
      ("1001001001010010", "01"), -- i=681
      ("1010001001010010", "10"), -- i=682
      ("1011001001010010", "11"), -- i=683
      ("1000001001010011", "00"), -- i=684
      ("1001001001010011", "01"), -- i=685
      ("1010001001010011", "10"), -- i=686
      ("1011001001010011", "11"), -- i=687
      ("1000001001010100", "00"), -- i=688
      ("1001001001010100", "01"), -- i=689
      ("1010001001010100", "10"), -- i=690
      ("1011001001010100", "11"), -- i=691
      ("1000001001010101", "00"), -- i=692
      ("1001001001010101", "01"), -- i=693
      ("1010001001010101", "10"), -- i=694
      ("1011001001010101", "11"), -- i=695
      ("1000001001010110", "00"), -- i=696
      ("1001001001010110", "01"), -- i=697
      ("1010001001010110", "10"), -- i=698
      ("1011001001010110", "11"), -- i=699
      ("1000001001010111", "00"), -- i=700
      ("1001001001010111", "01"), -- i=701
      ("1010001001010111", "10"), -- i=702
      ("1011001001010111", "11"), -- i=703
      ("1000001001100000", "00"), -- i=704
      ("1001001001100000", "01"), -- i=705
      ("1010001001100000", "10"), -- i=706
      ("1011001001100000", "11"), -- i=707
      ("1000001001100001", "00"), -- i=708
      ("1001001001100001", "01"), -- i=709
      ("1010001001100001", "10"), -- i=710
      ("1011001001100001", "11"), -- i=711
      ("1000001001100010", "00"), -- i=712
      ("1001001001100010", "01"), -- i=713
      ("1010001001100010", "10"), -- i=714
      ("1011001001100010", "11"), -- i=715
      ("1000001001100011", "00"), -- i=716
      ("1001001001100011", "01"), -- i=717
      ("1010001001100011", "10"), -- i=718
      ("1011001001100011", "11"), -- i=719
      ("1000001001100100", "00"), -- i=720
      ("1001001001100100", "01"), -- i=721
      ("1010001001100100", "10"), -- i=722
      ("1011001001100100", "11"), -- i=723
      ("1000001001100101", "00"), -- i=724
      ("1001001001100101", "01"), -- i=725
      ("1010001001100101", "10"), -- i=726
      ("1011001001100101", "11"), -- i=727
      ("1000001001100110", "00"), -- i=728
      ("1001001001100110", "01"), -- i=729
      ("1010001001100110", "10"), -- i=730
      ("1011001001100110", "11"), -- i=731
      ("1000001001100111", "00"), -- i=732
      ("1001001001100111", "01"), -- i=733
      ("1010001001100111", "10"), -- i=734
      ("1011001001100111", "11"), -- i=735
      ("1000001001110000", "00"), -- i=736
      ("1001001001110000", "01"), -- i=737
      ("1010001001110000", "10"), -- i=738
      ("1011001001110000", "11"), -- i=739
      ("1000001001110001", "00"), -- i=740
      ("1001001001110001", "01"), -- i=741
      ("1010001001110001", "10"), -- i=742
      ("1011001001110001", "11"), -- i=743
      ("1000001001110010", "00"), -- i=744
      ("1001001001110010", "01"), -- i=745
      ("1010001001110010", "10"), -- i=746
      ("1011001001110010", "11"), -- i=747
      ("1000001001110011", "00"), -- i=748
      ("1001001001110011", "01"), -- i=749
      ("1010001001110011", "10"), -- i=750
      ("1011001001110011", "11"), -- i=751
      ("1000001001110100", "00"), -- i=752
      ("1001001001110100", "01"), -- i=753
      ("1010001001110100", "10"), -- i=754
      ("1011001001110100", "11"), -- i=755
      ("1000001001110101", "00"), -- i=756
      ("1001001001110101", "01"), -- i=757
      ("1010001001110101", "10"), -- i=758
      ("1011001001110101", "11"), -- i=759
      ("1000001001110110", "00"), -- i=760
      ("1001001001110110", "01"), -- i=761
      ("1010001001110110", "10"), -- i=762
      ("1011001001110110", "11"), -- i=763
      ("1000001001110111", "00"), -- i=764
      ("1001001001110111", "01"), -- i=765
      ("1010001001110111", "10"), -- i=766
      ("1011001001110111", "11"), -- i=767
      ("1000001100000000", "00"), -- i=768
      ("1001001100000000", "01"), -- i=769
      ("1010001100000000", "10"), -- i=770
      ("1011001100000000", "11"), -- i=771
      ("1000001100000001", "00"), -- i=772
      ("1001001100000001", "01"), -- i=773
      ("1010001100000001", "10"), -- i=774
      ("1011001100000001", "11"), -- i=775
      ("1000001100000010", "00"), -- i=776
      ("1001001100000010", "01"), -- i=777
      ("1010001100000010", "10"), -- i=778
      ("1011001100000010", "11"), -- i=779
      ("1000001100000011", "00"), -- i=780
      ("1001001100000011", "01"), -- i=781
      ("1010001100000011", "10"), -- i=782
      ("1011001100000011", "11"), -- i=783
      ("1000001100000100", "00"), -- i=784
      ("1001001100000100", "01"), -- i=785
      ("1010001100000100", "10"), -- i=786
      ("1011001100000100", "11"), -- i=787
      ("1000001100000101", "00"), -- i=788
      ("1001001100000101", "01"), -- i=789
      ("1010001100000101", "10"), -- i=790
      ("1011001100000101", "11"), -- i=791
      ("1000001100000110", "00"), -- i=792
      ("1001001100000110", "01"), -- i=793
      ("1010001100000110", "10"), -- i=794
      ("1011001100000110", "11"), -- i=795
      ("1000001100000111", "00"), -- i=796
      ("1001001100000111", "01"), -- i=797
      ("1010001100000111", "10"), -- i=798
      ("1011001100000111", "11"), -- i=799
      ("1000001100010000", "00"), -- i=800
      ("1001001100010000", "01"), -- i=801
      ("1010001100010000", "10"), -- i=802
      ("1011001100010000", "11"), -- i=803
      ("1000001100010001", "00"), -- i=804
      ("1001001100010001", "01"), -- i=805
      ("1010001100010001", "10"), -- i=806
      ("1011001100010001", "11"), -- i=807
      ("1000001100010010", "00"), -- i=808
      ("1001001100010010", "01"), -- i=809
      ("1010001100010010", "10"), -- i=810
      ("1011001100010010", "11"), -- i=811
      ("1000001100010011", "00"), -- i=812
      ("1001001100010011", "01"), -- i=813
      ("1010001100010011", "10"), -- i=814
      ("1011001100010011", "11"), -- i=815
      ("1000001100010100", "00"), -- i=816
      ("1001001100010100", "01"), -- i=817
      ("1010001100010100", "10"), -- i=818
      ("1011001100010100", "11"), -- i=819
      ("1000001100010101", "00"), -- i=820
      ("1001001100010101", "01"), -- i=821
      ("1010001100010101", "10"), -- i=822
      ("1011001100010101", "11"), -- i=823
      ("1000001100010110", "00"), -- i=824
      ("1001001100010110", "01"), -- i=825
      ("1010001100010110", "10"), -- i=826
      ("1011001100010110", "11"), -- i=827
      ("1000001100010111", "00"), -- i=828
      ("1001001100010111", "01"), -- i=829
      ("1010001100010111", "10"), -- i=830
      ("1011001100010111", "11"), -- i=831
      ("1000001100100000", "00"), -- i=832
      ("1001001100100000", "01"), -- i=833
      ("1010001100100000", "10"), -- i=834
      ("1011001100100000", "11"), -- i=835
      ("1000001100100001", "00"), -- i=836
      ("1001001100100001", "01"), -- i=837
      ("1010001100100001", "10"), -- i=838
      ("1011001100100001", "11"), -- i=839
      ("1000001100100010", "00"), -- i=840
      ("1001001100100010", "01"), -- i=841
      ("1010001100100010", "10"), -- i=842
      ("1011001100100010", "11"), -- i=843
      ("1000001100100011", "00"), -- i=844
      ("1001001100100011", "01"), -- i=845
      ("1010001100100011", "10"), -- i=846
      ("1011001100100011", "11"), -- i=847
      ("1000001100100100", "00"), -- i=848
      ("1001001100100100", "01"), -- i=849
      ("1010001100100100", "10"), -- i=850
      ("1011001100100100", "11"), -- i=851
      ("1000001100100101", "00"), -- i=852
      ("1001001100100101", "01"), -- i=853
      ("1010001100100101", "10"), -- i=854
      ("1011001100100101", "11"), -- i=855
      ("1000001100100110", "00"), -- i=856
      ("1001001100100110", "01"), -- i=857
      ("1010001100100110", "10"), -- i=858
      ("1011001100100110", "11"), -- i=859
      ("1000001100100111", "00"), -- i=860
      ("1001001100100111", "01"), -- i=861
      ("1010001100100111", "10"), -- i=862
      ("1011001100100111", "11"), -- i=863
      ("1000001100110000", "00"), -- i=864
      ("1001001100110000", "01"), -- i=865
      ("1010001100110000", "10"), -- i=866
      ("1011001100110000", "11"), -- i=867
      ("1000001100110001", "00"), -- i=868
      ("1001001100110001", "01"), -- i=869
      ("1010001100110001", "10"), -- i=870
      ("1011001100110001", "11"), -- i=871
      ("1000001100110010", "00"), -- i=872
      ("1001001100110010", "01"), -- i=873
      ("1010001100110010", "10"), -- i=874
      ("1011001100110010", "11"), -- i=875
      ("1000001100110011", "00"), -- i=876
      ("1001001100110011", "01"), -- i=877
      ("1010001100110011", "10"), -- i=878
      ("1011001100110011", "11"), -- i=879
      ("1000001100110100", "00"), -- i=880
      ("1001001100110100", "01"), -- i=881
      ("1010001100110100", "10"), -- i=882
      ("1011001100110100", "11"), -- i=883
      ("1000001100110101", "00"), -- i=884
      ("1001001100110101", "01"), -- i=885
      ("1010001100110101", "10"), -- i=886
      ("1011001100110101", "11"), -- i=887
      ("1000001100110110", "00"), -- i=888
      ("1001001100110110", "01"), -- i=889
      ("1010001100110110", "10"), -- i=890
      ("1011001100110110", "11"), -- i=891
      ("1000001100110111", "00"), -- i=892
      ("1001001100110111", "01"), -- i=893
      ("1010001100110111", "10"), -- i=894
      ("1011001100110111", "11"), -- i=895
      ("1000001101000000", "00"), -- i=896
      ("1001001101000000", "01"), -- i=897
      ("1010001101000000", "10"), -- i=898
      ("1011001101000000", "11"), -- i=899
      ("1000001101000001", "00"), -- i=900
      ("1001001101000001", "01"), -- i=901
      ("1010001101000001", "10"), -- i=902
      ("1011001101000001", "11"), -- i=903
      ("1000001101000010", "00"), -- i=904
      ("1001001101000010", "01"), -- i=905
      ("1010001101000010", "10"), -- i=906
      ("1011001101000010", "11"), -- i=907
      ("1000001101000011", "00"), -- i=908
      ("1001001101000011", "01"), -- i=909
      ("1010001101000011", "10"), -- i=910
      ("1011001101000011", "11"), -- i=911
      ("1000001101000100", "00"), -- i=912
      ("1001001101000100", "01"), -- i=913
      ("1010001101000100", "10"), -- i=914
      ("1011001101000100", "11"), -- i=915
      ("1000001101000101", "00"), -- i=916
      ("1001001101000101", "01"), -- i=917
      ("1010001101000101", "10"), -- i=918
      ("1011001101000101", "11"), -- i=919
      ("1000001101000110", "00"), -- i=920
      ("1001001101000110", "01"), -- i=921
      ("1010001101000110", "10"), -- i=922
      ("1011001101000110", "11"), -- i=923
      ("1000001101000111", "00"), -- i=924
      ("1001001101000111", "01"), -- i=925
      ("1010001101000111", "10"), -- i=926
      ("1011001101000111", "11"), -- i=927
      ("1000001101010000", "00"), -- i=928
      ("1001001101010000", "01"), -- i=929
      ("1010001101010000", "10"), -- i=930
      ("1011001101010000", "11"), -- i=931
      ("1000001101010001", "00"), -- i=932
      ("1001001101010001", "01"), -- i=933
      ("1010001101010001", "10"), -- i=934
      ("1011001101010001", "11"), -- i=935
      ("1000001101010010", "00"), -- i=936
      ("1001001101010010", "01"), -- i=937
      ("1010001101010010", "10"), -- i=938
      ("1011001101010010", "11"), -- i=939
      ("1000001101010011", "00"), -- i=940
      ("1001001101010011", "01"), -- i=941
      ("1010001101010011", "10"), -- i=942
      ("1011001101010011", "11"), -- i=943
      ("1000001101010100", "00"), -- i=944
      ("1001001101010100", "01"), -- i=945
      ("1010001101010100", "10"), -- i=946
      ("1011001101010100", "11"), -- i=947
      ("1000001101010101", "00"), -- i=948
      ("1001001101010101", "01"), -- i=949
      ("1010001101010101", "10"), -- i=950
      ("1011001101010101", "11"), -- i=951
      ("1000001101010110", "00"), -- i=952
      ("1001001101010110", "01"), -- i=953
      ("1010001101010110", "10"), -- i=954
      ("1011001101010110", "11"), -- i=955
      ("1000001101010111", "00"), -- i=956
      ("1001001101010111", "01"), -- i=957
      ("1010001101010111", "10"), -- i=958
      ("1011001101010111", "11"), -- i=959
      ("1000001101100000", "00"), -- i=960
      ("1001001101100000", "01"), -- i=961
      ("1010001101100000", "10"), -- i=962
      ("1011001101100000", "11"), -- i=963
      ("1000001101100001", "00"), -- i=964
      ("1001001101100001", "01"), -- i=965
      ("1010001101100001", "10"), -- i=966
      ("1011001101100001", "11"), -- i=967
      ("1000001101100010", "00"), -- i=968
      ("1001001101100010", "01"), -- i=969
      ("1010001101100010", "10"), -- i=970
      ("1011001101100010", "11"), -- i=971
      ("1000001101100011", "00"), -- i=972
      ("1001001101100011", "01"), -- i=973
      ("1010001101100011", "10"), -- i=974
      ("1011001101100011", "11"), -- i=975
      ("1000001101100100", "00"), -- i=976
      ("1001001101100100", "01"), -- i=977
      ("1010001101100100", "10"), -- i=978
      ("1011001101100100", "11"), -- i=979
      ("1000001101100101", "00"), -- i=980
      ("1001001101100101", "01"), -- i=981
      ("1010001101100101", "10"), -- i=982
      ("1011001101100101", "11"), -- i=983
      ("1000001101100110", "00"), -- i=984
      ("1001001101100110", "01"), -- i=985
      ("1010001101100110", "10"), -- i=986
      ("1011001101100110", "11"), -- i=987
      ("1000001101100111", "00"), -- i=988
      ("1001001101100111", "01"), -- i=989
      ("1010001101100111", "10"), -- i=990
      ("1011001101100111", "11"), -- i=991
      ("1000001101110000", "00"), -- i=992
      ("1001001101110000", "01"), -- i=993
      ("1010001101110000", "10"), -- i=994
      ("1011001101110000", "11"), -- i=995
      ("1000001101110001", "00"), -- i=996
      ("1001001101110001", "01"), -- i=997
      ("1010001101110001", "10"), -- i=998
      ("1011001101110001", "11"), -- i=999
      ("1000001101110010", "00"), -- i=1000
      ("1001001101110010", "01"), -- i=1001
      ("1010001101110010", "10"), -- i=1002
      ("1011001101110010", "11"), -- i=1003
      ("1000001101110011", "00"), -- i=1004
      ("1001001101110011", "01"), -- i=1005
      ("1010001101110011", "10"), -- i=1006
      ("1011001101110011", "11"), -- i=1007
      ("1000001101110100", "00"), -- i=1008
      ("1001001101110100", "01"), -- i=1009
      ("1010001101110100", "10"), -- i=1010
      ("1011001101110100", "11"), -- i=1011
      ("1000001101110101", "00"), -- i=1012
      ("1001001101110101", "01"), -- i=1013
      ("1010001101110101", "10"), -- i=1014
      ("1011001101110101", "11"), -- i=1015
      ("1000001101110110", "00"), -- i=1016
      ("1001001101110110", "01"), -- i=1017
      ("1010001101110110", "10"), -- i=1018
      ("1011001101110110", "11"), -- i=1019
      ("1000001101110111", "00"), -- i=1020
      ("1001001101110111", "01"), -- i=1021
      ("1010001101110111", "10"), -- i=1022
      ("1011001101110111", "11"), -- i=1023
      ("1000010000000000", "00"), -- i=1024
      ("1001010000000000", "01"), -- i=1025
      ("1010010000000000", "10"), -- i=1026
      ("1011010000000000", "11"), -- i=1027
      ("1000010000000001", "00"), -- i=1028
      ("1001010000000001", "01"), -- i=1029
      ("1010010000000001", "10"), -- i=1030
      ("1011010000000001", "11"), -- i=1031
      ("1000010000000010", "00"), -- i=1032
      ("1001010000000010", "01"), -- i=1033
      ("1010010000000010", "10"), -- i=1034
      ("1011010000000010", "11"), -- i=1035
      ("1000010000000011", "00"), -- i=1036
      ("1001010000000011", "01"), -- i=1037
      ("1010010000000011", "10"), -- i=1038
      ("1011010000000011", "11"), -- i=1039
      ("1000010000000100", "00"), -- i=1040
      ("1001010000000100", "01"), -- i=1041
      ("1010010000000100", "10"), -- i=1042
      ("1011010000000100", "11"), -- i=1043
      ("1000010000000101", "00"), -- i=1044
      ("1001010000000101", "01"), -- i=1045
      ("1010010000000101", "10"), -- i=1046
      ("1011010000000101", "11"), -- i=1047
      ("1000010000000110", "00"), -- i=1048
      ("1001010000000110", "01"), -- i=1049
      ("1010010000000110", "10"), -- i=1050
      ("1011010000000110", "11"), -- i=1051
      ("1000010000000111", "00"), -- i=1052
      ("1001010000000111", "01"), -- i=1053
      ("1010010000000111", "10"), -- i=1054
      ("1011010000000111", "11"), -- i=1055
      ("1000010000010000", "00"), -- i=1056
      ("1001010000010000", "01"), -- i=1057
      ("1010010000010000", "10"), -- i=1058
      ("1011010000010000", "11"), -- i=1059
      ("1000010000010001", "00"), -- i=1060
      ("1001010000010001", "01"), -- i=1061
      ("1010010000010001", "10"), -- i=1062
      ("1011010000010001", "11"), -- i=1063
      ("1000010000010010", "00"), -- i=1064
      ("1001010000010010", "01"), -- i=1065
      ("1010010000010010", "10"), -- i=1066
      ("1011010000010010", "11"), -- i=1067
      ("1000010000010011", "00"), -- i=1068
      ("1001010000010011", "01"), -- i=1069
      ("1010010000010011", "10"), -- i=1070
      ("1011010000010011", "11"), -- i=1071
      ("1000010000010100", "00"), -- i=1072
      ("1001010000010100", "01"), -- i=1073
      ("1010010000010100", "10"), -- i=1074
      ("1011010000010100", "11"), -- i=1075
      ("1000010000010101", "00"), -- i=1076
      ("1001010000010101", "01"), -- i=1077
      ("1010010000010101", "10"), -- i=1078
      ("1011010000010101", "11"), -- i=1079
      ("1000010000010110", "00"), -- i=1080
      ("1001010000010110", "01"), -- i=1081
      ("1010010000010110", "10"), -- i=1082
      ("1011010000010110", "11"), -- i=1083
      ("1000010000010111", "00"), -- i=1084
      ("1001010000010111", "01"), -- i=1085
      ("1010010000010111", "10"), -- i=1086
      ("1011010000010111", "11"), -- i=1087
      ("1000010000100000", "00"), -- i=1088
      ("1001010000100000", "01"), -- i=1089
      ("1010010000100000", "10"), -- i=1090
      ("1011010000100000", "11"), -- i=1091
      ("1000010000100001", "00"), -- i=1092
      ("1001010000100001", "01"), -- i=1093
      ("1010010000100001", "10"), -- i=1094
      ("1011010000100001", "11"), -- i=1095
      ("1000010000100010", "00"), -- i=1096
      ("1001010000100010", "01"), -- i=1097
      ("1010010000100010", "10"), -- i=1098
      ("1011010000100010", "11"), -- i=1099
      ("1000010000100011", "00"), -- i=1100
      ("1001010000100011", "01"), -- i=1101
      ("1010010000100011", "10"), -- i=1102
      ("1011010000100011", "11"), -- i=1103
      ("1000010000100100", "00"), -- i=1104
      ("1001010000100100", "01"), -- i=1105
      ("1010010000100100", "10"), -- i=1106
      ("1011010000100100", "11"), -- i=1107
      ("1000010000100101", "00"), -- i=1108
      ("1001010000100101", "01"), -- i=1109
      ("1010010000100101", "10"), -- i=1110
      ("1011010000100101", "11"), -- i=1111
      ("1000010000100110", "00"), -- i=1112
      ("1001010000100110", "01"), -- i=1113
      ("1010010000100110", "10"), -- i=1114
      ("1011010000100110", "11"), -- i=1115
      ("1000010000100111", "00"), -- i=1116
      ("1001010000100111", "01"), -- i=1117
      ("1010010000100111", "10"), -- i=1118
      ("1011010000100111", "11"), -- i=1119
      ("1000010000110000", "00"), -- i=1120
      ("1001010000110000", "01"), -- i=1121
      ("1010010000110000", "10"), -- i=1122
      ("1011010000110000", "11"), -- i=1123
      ("1000010000110001", "00"), -- i=1124
      ("1001010000110001", "01"), -- i=1125
      ("1010010000110001", "10"), -- i=1126
      ("1011010000110001", "11"), -- i=1127
      ("1000010000110010", "00"), -- i=1128
      ("1001010000110010", "01"), -- i=1129
      ("1010010000110010", "10"), -- i=1130
      ("1011010000110010", "11"), -- i=1131
      ("1000010000110011", "00"), -- i=1132
      ("1001010000110011", "01"), -- i=1133
      ("1010010000110011", "10"), -- i=1134
      ("1011010000110011", "11"), -- i=1135
      ("1000010000110100", "00"), -- i=1136
      ("1001010000110100", "01"), -- i=1137
      ("1010010000110100", "10"), -- i=1138
      ("1011010000110100", "11"), -- i=1139
      ("1000010000110101", "00"), -- i=1140
      ("1001010000110101", "01"), -- i=1141
      ("1010010000110101", "10"), -- i=1142
      ("1011010000110101", "11"), -- i=1143
      ("1000010000110110", "00"), -- i=1144
      ("1001010000110110", "01"), -- i=1145
      ("1010010000110110", "10"), -- i=1146
      ("1011010000110110", "11"), -- i=1147
      ("1000010000110111", "00"), -- i=1148
      ("1001010000110111", "01"), -- i=1149
      ("1010010000110111", "10"), -- i=1150
      ("1011010000110111", "11"), -- i=1151
      ("1000010001000000", "00"), -- i=1152
      ("1001010001000000", "01"), -- i=1153
      ("1010010001000000", "10"), -- i=1154
      ("1011010001000000", "11"), -- i=1155
      ("1000010001000001", "00"), -- i=1156
      ("1001010001000001", "01"), -- i=1157
      ("1010010001000001", "10"), -- i=1158
      ("1011010001000001", "11"), -- i=1159
      ("1000010001000010", "00"), -- i=1160
      ("1001010001000010", "01"), -- i=1161
      ("1010010001000010", "10"), -- i=1162
      ("1011010001000010", "11"), -- i=1163
      ("1000010001000011", "00"), -- i=1164
      ("1001010001000011", "01"), -- i=1165
      ("1010010001000011", "10"), -- i=1166
      ("1011010001000011", "11"), -- i=1167
      ("1000010001000100", "00"), -- i=1168
      ("1001010001000100", "01"), -- i=1169
      ("1010010001000100", "10"), -- i=1170
      ("1011010001000100", "11"), -- i=1171
      ("1000010001000101", "00"), -- i=1172
      ("1001010001000101", "01"), -- i=1173
      ("1010010001000101", "10"), -- i=1174
      ("1011010001000101", "11"), -- i=1175
      ("1000010001000110", "00"), -- i=1176
      ("1001010001000110", "01"), -- i=1177
      ("1010010001000110", "10"), -- i=1178
      ("1011010001000110", "11"), -- i=1179
      ("1000010001000111", "00"), -- i=1180
      ("1001010001000111", "01"), -- i=1181
      ("1010010001000111", "10"), -- i=1182
      ("1011010001000111", "11"), -- i=1183
      ("1000010001010000", "00"), -- i=1184
      ("1001010001010000", "01"), -- i=1185
      ("1010010001010000", "10"), -- i=1186
      ("1011010001010000", "11"), -- i=1187
      ("1000010001010001", "00"), -- i=1188
      ("1001010001010001", "01"), -- i=1189
      ("1010010001010001", "10"), -- i=1190
      ("1011010001010001", "11"), -- i=1191
      ("1000010001010010", "00"), -- i=1192
      ("1001010001010010", "01"), -- i=1193
      ("1010010001010010", "10"), -- i=1194
      ("1011010001010010", "11"), -- i=1195
      ("1000010001010011", "00"), -- i=1196
      ("1001010001010011", "01"), -- i=1197
      ("1010010001010011", "10"), -- i=1198
      ("1011010001010011", "11"), -- i=1199
      ("1000010001010100", "00"), -- i=1200
      ("1001010001010100", "01"), -- i=1201
      ("1010010001010100", "10"), -- i=1202
      ("1011010001010100", "11"), -- i=1203
      ("1000010001010101", "00"), -- i=1204
      ("1001010001010101", "01"), -- i=1205
      ("1010010001010101", "10"), -- i=1206
      ("1011010001010101", "11"), -- i=1207
      ("1000010001010110", "00"), -- i=1208
      ("1001010001010110", "01"), -- i=1209
      ("1010010001010110", "10"), -- i=1210
      ("1011010001010110", "11"), -- i=1211
      ("1000010001010111", "00"), -- i=1212
      ("1001010001010111", "01"), -- i=1213
      ("1010010001010111", "10"), -- i=1214
      ("1011010001010111", "11"), -- i=1215
      ("1000010001100000", "00"), -- i=1216
      ("1001010001100000", "01"), -- i=1217
      ("1010010001100000", "10"), -- i=1218
      ("1011010001100000", "11"), -- i=1219
      ("1000010001100001", "00"), -- i=1220
      ("1001010001100001", "01"), -- i=1221
      ("1010010001100001", "10"), -- i=1222
      ("1011010001100001", "11"), -- i=1223
      ("1000010001100010", "00"), -- i=1224
      ("1001010001100010", "01"), -- i=1225
      ("1010010001100010", "10"), -- i=1226
      ("1011010001100010", "11"), -- i=1227
      ("1000010001100011", "00"), -- i=1228
      ("1001010001100011", "01"), -- i=1229
      ("1010010001100011", "10"), -- i=1230
      ("1011010001100011", "11"), -- i=1231
      ("1000010001100100", "00"), -- i=1232
      ("1001010001100100", "01"), -- i=1233
      ("1010010001100100", "10"), -- i=1234
      ("1011010001100100", "11"), -- i=1235
      ("1000010001100101", "00"), -- i=1236
      ("1001010001100101", "01"), -- i=1237
      ("1010010001100101", "10"), -- i=1238
      ("1011010001100101", "11"), -- i=1239
      ("1000010001100110", "00"), -- i=1240
      ("1001010001100110", "01"), -- i=1241
      ("1010010001100110", "10"), -- i=1242
      ("1011010001100110", "11"), -- i=1243
      ("1000010001100111", "00"), -- i=1244
      ("1001010001100111", "01"), -- i=1245
      ("1010010001100111", "10"), -- i=1246
      ("1011010001100111", "11"), -- i=1247
      ("1000010001110000", "00"), -- i=1248
      ("1001010001110000", "01"), -- i=1249
      ("1010010001110000", "10"), -- i=1250
      ("1011010001110000", "11"), -- i=1251
      ("1000010001110001", "00"), -- i=1252
      ("1001010001110001", "01"), -- i=1253
      ("1010010001110001", "10"), -- i=1254
      ("1011010001110001", "11"), -- i=1255
      ("1000010001110010", "00"), -- i=1256
      ("1001010001110010", "01"), -- i=1257
      ("1010010001110010", "10"), -- i=1258
      ("1011010001110010", "11"), -- i=1259
      ("1000010001110011", "00"), -- i=1260
      ("1001010001110011", "01"), -- i=1261
      ("1010010001110011", "10"), -- i=1262
      ("1011010001110011", "11"), -- i=1263
      ("1000010001110100", "00"), -- i=1264
      ("1001010001110100", "01"), -- i=1265
      ("1010010001110100", "10"), -- i=1266
      ("1011010001110100", "11"), -- i=1267
      ("1000010001110101", "00"), -- i=1268
      ("1001010001110101", "01"), -- i=1269
      ("1010010001110101", "10"), -- i=1270
      ("1011010001110101", "11"), -- i=1271
      ("1000010001110110", "00"), -- i=1272
      ("1001010001110110", "01"), -- i=1273
      ("1010010001110110", "10"), -- i=1274
      ("1011010001110110", "11"), -- i=1275
      ("1000010001110111", "00"), -- i=1276
      ("1001010001110111", "01"), -- i=1277
      ("1010010001110111", "10"), -- i=1278
      ("1011010001110111", "11"), -- i=1279
      ("1000010100000000", "00"), -- i=1280
      ("1001010100000000", "01"), -- i=1281
      ("1010010100000000", "10"), -- i=1282
      ("1011010100000000", "11"), -- i=1283
      ("1000010100000001", "00"), -- i=1284
      ("1001010100000001", "01"), -- i=1285
      ("1010010100000001", "10"), -- i=1286
      ("1011010100000001", "11"), -- i=1287
      ("1000010100000010", "00"), -- i=1288
      ("1001010100000010", "01"), -- i=1289
      ("1010010100000010", "10"), -- i=1290
      ("1011010100000010", "11"), -- i=1291
      ("1000010100000011", "00"), -- i=1292
      ("1001010100000011", "01"), -- i=1293
      ("1010010100000011", "10"), -- i=1294
      ("1011010100000011", "11"), -- i=1295
      ("1000010100000100", "00"), -- i=1296
      ("1001010100000100", "01"), -- i=1297
      ("1010010100000100", "10"), -- i=1298
      ("1011010100000100", "11"), -- i=1299
      ("1000010100000101", "00"), -- i=1300
      ("1001010100000101", "01"), -- i=1301
      ("1010010100000101", "10"), -- i=1302
      ("1011010100000101", "11"), -- i=1303
      ("1000010100000110", "00"), -- i=1304
      ("1001010100000110", "01"), -- i=1305
      ("1010010100000110", "10"), -- i=1306
      ("1011010100000110", "11"), -- i=1307
      ("1000010100000111", "00"), -- i=1308
      ("1001010100000111", "01"), -- i=1309
      ("1010010100000111", "10"), -- i=1310
      ("1011010100000111", "11"), -- i=1311
      ("1000010100010000", "00"), -- i=1312
      ("1001010100010000", "01"), -- i=1313
      ("1010010100010000", "10"), -- i=1314
      ("1011010100010000", "11"), -- i=1315
      ("1000010100010001", "00"), -- i=1316
      ("1001010100010001", "01"), -- i=1317
      ("1010010100010001", "10"), -- i=1318
      ("1011010100010001", "11"), -- i=1319
      ("1000010100010010", "00"), -- i=1320
      ("1001010100010010", "01"), -- i=1321
      ("1010010100010010", "10"), -- i=1322
      ("1011010100010010", "11"), -- i=1323
      ("1000010100010011", "00"), -- i=1324
      ("1001010100010011", "01"), -- i=1325
      ("1010010100010011", "10"), -- i=1326
      ("1011010100010011", "11"), -- i=1327
      ("1000010100010100", "00"), -- i=1328
      ("1001010100010100", "01"), -- i=1329
      ("1010010100010100", "10"), -- i=1330
      ("1011010100010100", "11"), -- i=1331
      ("1000010100010101", "00"), -- i=1332
      ("1001010100010101", "01"), -- i=1333
      ("1010010100010101", "10"), -- i=1334
      ("1011010100010101", "11"), -- i=1335
      ("1000010100010110", "00"), -- i=1336
      ("1001010100010110", "01"), -- i=1337
      ("1010010100010110", "10"), -- i=1338
      ("1011010100010110", "11"), -- i=1339
      ("1000010100010111", "00"), -- i=1340
      ("1001010100010111", "01"), -- i=1341
      ("1010010100010111", "10"), -- i=1342
      ("1011010100010111", "11"), -- i=1343
      ("1000010100100000", "00"), -- i=1344
      ("1001010100100000", "01"), -- i=1345
      ("1010010100100000", "10"), -- i=1346
      ("1011010100100000", "11"), -- i=1347
      ("1000010100100001", "00"), -- i=1348
      ("1001010100100001", "01"), -- i=1349
      ("1010010100100001", "10"), -- i=1350
      ("1011010100100001", "11"), -- i=1351
      ("1000010100100010", "00"), -- i=1352
      ("1001010100100010", "01"), -- i=1353
      ("1010010100100010", "10"), -- i=1354
      ("1011010100100010", "11"), -- i=1355
      ("1000010100100011", "00"), -- i=1356
      ("1001010100100011", "01"), -- i=1357
      ("1010010100100011", "10"), -- i=1358
      ("1011010100100011", "11"), -- i=1359
      ("1000010100100100", "00"), -- i=1360
      ("1001010100100100", "01"), -- i=1361
      ("1010010100100100", "10"), -- i=1362
      ("1011010100100100", "11"), -- i=1363
      ("1000010100100101", "00"), -- i=1364
      ("1001010100100101", "01"), -- i=1365
      ("1010010100100101", "10"), -- i=1366
      ("1011010100100101", "11"), -- i=1367
      ("1000010100100110", "00"), -- i=1368
      ("1001010100100110", "01"), -- i=1369
      ("1010010100100110", "10"), -- i=1370
      ("1011010100100110", "11"), -- i=1371
      ("1000010100100111", "00"), -- i=1372
      ("1001010100100111", "01"), -- i=1373
      ("1010010100100111", "10"), -- i=1374
      ("1011010100100111", "11"), -- i=1375
      ("1000010100110000", "00"), -- i=1376
      ("1001010100110000", "01"), -- i=1377
      ("1010010100110000", "10"), -- i=1378
      ("1011010100110000", "11"), -- i=1379
      ("1000010100110001", "00"), -- i=1380
      ("1001010100110001", "01"), -- i=1381
      ("1010010100110001", "10"), -- i=1382
      ("1011010100110001", "11"), -- i=1383
      ("1000010100110010", "00"), -- i=1384
      ("1001010100110010", "01"), -- i=1385
      ("1010010100110010", "10"), -- i=1386
      ("1011010100110010", "11"), -- i=1387
      ("1000010100110011", "00"), -- i=1388
      ("1001010100110011", "01"), -- i=1389
      ("1010010100110011", "10"), -- i=1390
      ("1011010100110011", "11"), -- i=1391
      ("1000010100110100", "00"), -- i=1392
      ("1001010100110100", "01"), -- i=1393
      ("1010010100110100", "10"), -- i=1394
      ("1011010100110100", "11"), -- i=1395
      ("1000010100110101", "00"), -- i=1396
      ("1001010100110101", "01"), -- i=1397
      ("1010010100110101", "10"), -- i=1398
      ("1011010100110101", "11"), -- i=1399
      ("1000010100110110", "00"), -- i=1400
      ("1001010100110110", "01"), -- i=1401
      ("1010010100110110", "10"), -- i=1402
      ("1011010100110110", "11"), -- i=1403
      ("1000010100110111", "00"), -- i=1404
      ("1001010100110111", "01"), -- i=1405
      ("1010010100110111", "10"), -- i=1406
      ("1011010100110111", "11"), -- i=1407
      ("1000010101000000", "00"), -- i=1408
      ("1001010101000000", "01"), -- i=1409
      ("1010010101000000", "10"), -- i=1410
      ("1011010101000000", "11"), -- i=1411
      ("1000010101000001", "00"), -- i=1412
      ("1001010101000001", "01"), -- i=1413
      ("1010010101000001", "10"), -- i=1414
      ("1011010101000001", "11"), -- i=1415
      ("1000010101000010", "00"), -- i=1416
      ("1001010101000010", "01"), -- i=1417
      ("1010010101000010", "10"), -- i=1418
      ("1011010101000010", "11"), -- i=1419
      ("1000010101000011", "00"), -- i=1420
      ("1001010101000011", "01"), -- i=1421
      ("1010010101000011", "10"), -- i=1422
      ("1011010101000011", "11"), -- i=1423
      ("1000010101000100", "00"), -- i=1424
      ("1001010101000100", "01"), -- i=1425
      ("1010010101000100", "10"), -- i=1426
      ("1011010101000100", "11"), -- i=1427
      ("1000010101000101", "00"), -- i=1428
      ("1001010101000101", "01"), -- i=1429
      ("1010010101000101", "10"), -- i=1430
      ("1011010101000101", "11"), -- i=1431
      ("1000010101000110", "00"), -- i=1432
      ("1001010101000110", "01"), -- i=1433
      ("1010010101000110", "10"), -- i=1434
      ("1011010101000110", "11"), -- i=1435
      ("1000010101000111", "00"), -- i=1436
      ("1001010101000111", "01"), -- i=1437
      ("1010010101000111", "10"), -- i=1438
      ("1011010101000111", "11"), -- i=1439
      ("1000010101010000", "00"), -- i=1440
      ("1001010101010000", "01"), -- i=1441
      ("1010010101010000", "10"), -- i=1442
      ("1011010101010000", "11"), -- i=1443
      ("1000010101010001", "00"), -- i=1444
      ("1001010101010001", "01"), -- i=1445
      ("1010010101010001", "10"), -- i=1446
      ("1011010101010001", "11"), -- i=1447
      ("1000010101010010", "00"), -- i=1448
      ("1001010101010010", "01"), -- i=1449
      ("1010010101010010", "10"), -- i=1450
      ("1011010101010010", "11"), -- i=1451
      ("1000010101010011", "00"), -- i=1452
      ("1001010101010011", "01"), -- i=1453
      ("1010010101010011", "10"), -- i=1454
      ("1011010101010011", "11"), -- i=1455
      ("1000010101010100", "00"), -- i=1456
      ("1001010101010100", "01"), -- i=1457
      ("1010010101010100", "10"), -- i=1458
      ("1011010101010100", "11"), -- i=1459
      ("1000010101010101", "00"), -- i=1460
      ("1001010101010101", "01"), -- i=1461
      ("1010010101010101", "10"), -- i=1462
      ("1011010101010101", "11"), -- i=1463
      ("1000010101010110", "00"), -- i=1464
      ("1001010101010110", "01"), -- i=1465
      ("1010010101010110", "10"), -- i=1466
      ("1011010101010110", "11"), -- i=1467
      ("1000010101010111", "00"), -- i=1468
      ("1001010101010111", "01"), -- i=1469
      ("1010010101010111", "10"), -- i=1470
      ("1011010101010111", "11"), -- i=1471
      ("1000010101100000", "00"), -- i=1472
      ("1001010101100000", "01"), -- i=1473
      ("1010010101100000", "10"), -- i=1474
      ("1011010101100000", "11"), -- i=1475
      ("1000010101100001", "00"), -- i=1476
      ("1001010101100001", "01"), -- i=1477
      ("1010010101100001", "10"), -- i=1478
      ("1011010101100001", "11"), -- i=1479
      ("1000010101100010", "00"), -- i=1480
      ("1001010101100010", "01"), -- i=1481
      ("1010010101100010", "10"), -- i=1482
      ("1011010101100010", "11"), -- i=1483
      ("1000010101100011", "00"), -- i=1484
      ("1001010101100011", "01"), -- i=1485
      ("1010010101100011", "10"), -- i=1486
      ("1011010101100011", "11"), -- i=1487
      ("1000010101100100", "00"), -- i=1488
      ("1001010101100100", "01"), -- i=1489
      ("1010010101100100", "10"), -- i=1490
      ("1011010101100100", "11"), -- i=1491
      ("1000010101100101", "00"), -- i=1492
      ("1001010101100101", "01"), -- i=1493
      ("1010010101100101", "10"), -- i=1494
      ("1011010101100101", "11"), -- i=1495
      ("1000010101100110", "00"), -- i=1496
      ("1001010101100110", "01"), -- i=1497
      ("1010010101100110", "10"), -- i=1498
      ("1011010101100110", "11"), -- i=1499
      ("1000010101100111", "00"), -- i=1500
      ("1001010101100111", "01"), -- i=1501
      ("1010010101100111", "10"), -- i=1502
      ("1011010101100111", "11"), -- i=1503
      ("1000010101110000", "00"), -- i=1504
      ("1001010101110000", "01"), -- i=1505
      ("1010010101110000", "10"), -- i=1506
      ("1011010101110000", "11"), -- i=1507
      ("1000010101110001", "00"), -- i=1508
      ("1001010101110001", "01"), -- i=1509
      ("1010010101110001", "10"), -- i=1510
      ("1011010101110001", "11"), -- i=1511
      ("1000010101110010", "00"), -- i=1512
      ("1001010101110010", "01"), -- i=1513
      ("1010010101110010", "10"), -- i=1514
      ("1011010101110010", "11"), -- i=1515
      ("1000010101110011", "00"), -- i=1516
      ("1001010101110011", "01"), -- i=1517
      ("1010010101110011", "10"), -- i=1518
      ("1011010101110011", "11"), -- i=1519
      ("1000010101110100", "00"), -- i=1520
      ("1001010101110100", "01"), -- i=1521
      ("1010010101110100", "10"), -- i=1522
      ("1011010101110100", "11"), -- i=1523
      ("1000010101110101", "00"), -- i=1524
      ("1001010101110101", "01"), -- i=1525
      ("1010010101110101", "10"), -- i=1526
      ("1011010101110101", "11"), -- i=1527
      ("1000010101110110", "00"), -- i=1528
      ("1001010101110110", "01"), -- i=1529
      ("1010010101110110", "10"), -- i=1530
      ("1011010101110110", "11"), -- i=1531
      ("1000010101110111", "00"), -- i=1532
      ("1001010101110111", "01"), -- i=1533
      ("1010010101110111", "10"), -- i=1534
      ("1011010101110111", "11"), -- i=1535
      ("1000011000000000", "00"), -- i=1536
      ("1001011000000000", "01"), -- i=1537
      ("1010011000000000", "10"), -- i=1538
      ("1011011000000000", "11"), -- i=1539
      ("1000011000000001", "00"), -- i=1540
      ("1001011000000001", "01"), -- i=1541
      ("1010011000000001", "10"), -- i=1542
      ("1011011000000001", "11"), -- i=1543
      ("1000011000000010", "00"), -- i=1544
      ("1001011000000010", "01"), -- i=1545
      ("1010011000000010", "10"), -- i=1546
      ("1011011000000010", "11"), -- i=1547
      ("1000011000000011", "00"), -- i=1548
      ("1001011000000011", "01"), -- i=1549
      ("1010011000000011", "10"), -- i=1550
      ("1011011000000011", "11"), -- i=1551
      ("1000011000000100", "00"), -- i=1552
      ("1001011000000100", "01"), -- i=1553
      ("1010011000000100", "10"), -- i=1554
      ("1011011000000100", "11"), -- i=1555
      ("1000011000000101", "00"), -- i=1556
      ("1001011000000101", "01"), -- i=1557
      ("1010011000000101", "10"), -- i=1558
      ("1011011000000101", "11"), -- i=1559
      ("1000011000000110", "00"), -- i=1560
      ("1001011000000110", "01"), -- i=1561
      ("1010011000000110", "10"), -- i=1562
      ("1011011000000110", "11"), -- i=1563
      ("1000011000000111", "00"), -- i=1564
      ("1001011000000111", "01"), -- i=1565
      ("1010011000000111", "10"), -- i=1566
      ("1011011000000111", "11"), -- i=1567
      ("1000011000010000", "00"), -- i=1568
      ("1001011000010000", "01"), -- i=1569
      ("1010011000010000", "10"), -- i=1570
      ("1011011000010000", "11"), -- i=1571
      ("1000011000010001", "00"), -- i=1572
      ("1001011000010001", "01"), -- i=1573
      ("1010011000010001", "10"), -- i=1574
      ("1011011000010001", "11"), -- i=1575
      ("1000011000010010", "00"), -- i=1576
      ("1001011000010010", "01"), -- i=1577
      ("1010011000010010", "10"), -- i=1578
      ("1011011000010010", "11"), -- i=1579
      ("1000011000010011", "00"), -- i=1580
      ("1001011000010011", "01"), -- i=1581
      ("1010011000010011", "10"), -- i=1582
      ("1011011000010011", "11"), -- i=1583
      ("1000011000010100", "00"), -- i=1584
      ("1001011000010100", "01"), -- i=1585
      ("1010011000010100", "10"), -- i=1586
      ("1011011000010100", "11"), -- i=1587
      ("1000011000010101", "00"), -- i=1588
      ("1001011000010101", "01"), -- i=1589
      ("1010011000010101", "10"), -- i=1590
      ("1011011000010101", "11"), -- i=1591
      ("1000011000010110", "00"), -- i=1592
      ("1001011000010110", "01"), -- i=1593
      ("1010011000010110", "10"), -- i=1594
      ("1011011000010110", "11"), -- i=1595
      ("1000011000010111", "00"), -- i=1596
      ("1001011000010111", "01"), -- i=1597
      ("1010011000010111", "10"), -- i=1598
      ("1011011000010111", "11"), -- i=1599
      ("1000011000100000", "00"), -- i=1600
      ("1001011000100000", "01"), -- i=1601
      ("1010011000100000", "10"), -- i=1602
      ("1011011000100000", "11"), -- i=1603
      ("1000011000100001", "00"), -- i=1604
      ("1001011000100001", "01"), -- i=1605
      ("1010011000100001", "10"), -- i=1606
      ("1011011000100001", "11"), -- i=1607
      ("1000011000100010", "00"), -- i=1608
      ("1001011000100010", "01"), -- i=1609
      ("1010011000100010", "10"), -- i=1610
      ("1011011000100010", "11"), -- i=1611
      ("1000011000100011", "00"), -- i=1612
      ("1001011000100011", "01"), -- i=1613
      ("1010011000100011", "10"), -- i=1614
      ("1011011000100011", "11"), -- i=1615
      ("1000011000100100", "00"), -- i=1616
      ("1001011000100100", "01"), -- i=1617
      ("1010011000100100", "10"), -- i=1618
      ("1011011000100100", "11"), -- i=1619
      ("1000011000100101", "00"), -- i=1620
      ("1001011000100101", "01"), -- i=1621
      ("1010011000100101", "10"), -- i=1622
      ("1011011000100101", "11"), -- i=1623
      ("1000011000100110", "00"), -- i=1624
      ("1001011000100110", "01"), -- i=1625
      ("1010011000100110", "10"), -- i=1626
      ("1011011000100110", "11"), -- i=1627
      ("1000011000100111", "00"), -- i=1628
      ("1001011000100111", "01"), -- i=1629
      ("1010011000100111", "10"), -- i=1630
      ("1011011000100111", "11"), -- i=1631
      ("1000011000110000", "00"), -- i=1632
      ("1001011000110000", "01"), -- i=1633
      ("1010011000110000", "10"), -- i=1634
      ("1011011000110000", "11"), -- i=1635
      ("1000011000110001", "00"), -- i=1636
      ("1001011000110001", "01"), -- i=1637
      ("1010011000110001", "10"), -- i=1638
      ("1011011000110001", "11"), -- i=1639
      ("1000011000110010", "00"), -- i=1640
      ("1001011000110010", "01"), -- i=1641
      ("1010011000110010", "10"), -- i=1642
      ("1011011000110010", "11"), -- i=1643
      ("1000011000110011", "00"), -- i=1644
      ("1001011000110011", "01"), -- i=1645
      ("1010011000110011", "10"), -- i=1646
      ("1011011000110011", "11"), -- i=1647
      ("1000011000110100", "00"), -- i=1648
      ("1001011000110100", "01"), -- i=1649
      ("1010011000110100", "10"), -- i=1650
      ("1011011000110100", "11"), -- i=1651
      ("1000011000110101", "00"), -- i=1652
      ("1001011000110101", "01"), -- i=1653
      ("1010011000110101", "10"), -- i=1654
      ("1011011000110101", "11"), -- i=1655
      ("1000011000110110", "00"), -- i=1656
      ("1001011000110110", "01"), -- i=1657
      ("1010011000110110", "10"), -- i=1658
      ("1011011000110110", "11"), -- i=1659
      ("1000011000110111", "00"), -- i=1660
      ("1001011000110111", "01"), -- i=1661
      ("1010011000110111", "10"), -- i=1662
      ("1011011000110111", "11"), -- i=1663
      ("1000011001000000", "00"), -- i=1664
      ("1001011001000000", "01"), -- i=1665
      ("1010011001000000", "10"), -- i=1666
      ("1011011001000000", "11"), -- i=1667
      ("1000011001000001", "00"), -- i=1668
      ("1001011001000001", "01"), -- i=1669
      ("1010011001000001", "10"), -- i=1670
      ("1011011001000001", "11"), -- i=1671
      ("1000011001000010", "00"), -- i=1672
      ("1001011001000010", "01"), -- i=1673
      ("1010011001000010", "10"), -- i=1674
      ("1011011001000010", "11"), -- i=1675
      ("1000011001000011", "00"), -- i=1676
      ("1001011001000011", "01"), -- i=1677
      ("1010011001000011", "10"), -- i=1678
      ("1011011001000011", "11"), -- i=1679
      ("1000011001000100", "00"), -- i=1680
      ("1001011001000100", "01"), -- i=1681
      ("1010011001000100", "10"), -- i=1682
      ("1011011001000100", "11"), -- i=1683
      ("1000011001000101", "00"), -- i=1684
      ("1001011001000101", "01"), -- i=1685
      ("1010011001000101", "10"), -- i=1686
      ("1011011001000101", "11"), -- i=1687
      ("1000011001000110", "00"), -- i=1688
      ("1001011001000110", "01"), -- i=1689
      ("1010011001000110", "10"), -- i=1690
      ("1011011001000110", "11"), -- i=1691
      ("1000011001000111", "00"), -- i=1692
      ("1001011001000111", "01"), -- i=1693
      ("1010011001000111", "10"), -- i=1694
      ("1011011001000111", "11"), -- i=1695
      ("1000011001010000", "00"), -- i=1696
      ("1001011001010000", "01"), -- i=1697
      ("1010011001010000", "10"), -- i=1698
      ("1011011001010000", "11"), -- i=1699
      ("1000011001010001", "00"), -- i=1700
      ("1001011001010001", "01"), -- i=1701
      ("1010011001010001", "10"), -- i=1702
      ("1011011001010001", "11"), -- i=1703
      ("1000011001010010", "00"), -- i=1704
      ("1001011001010010", "01"), -- i=1705
      ("1010011001010010", "10"), -- i=1706
      ("1011011001010010", "11"), -- i=1707
      ("1000011001010011", "00"), -- i=1708
      ("1001011001010011", "01"), -- i=1709
      ("1010011001010011", "10"), -- i=1710
      ("1011011001010011", "11"), -- i=1711
      ("1000011001010100", "00"), -- i=1712
      ("1001011001010100", "01"), -- i=1713
      ("1010011001010100", "10"), -- i=1714
      ("1011011001010100", "11"), -- i=1715
      ("1000011001010101", "00"), -- i=1716
      ("1001011001010101", "01"), -- i=1717
      ("1010011001010101", "10"), -- i=1718
      ("1011011001010101", "11"), -- i=1719
      ("1000011001010110", "00"), -- i=1720
      ("1001011001010110", "01"), -- i=1721
      ("1010011001010110", "10"), -- i=1722
      ("1011011001010110", "11"), -- i=1723
      ("1000011001010111", "00"), -- i=1724
      ("1001011001010111", "01"), -- i=1725
      ("1010011001010111", "10"), -- i=1726
      ("1011011001010111", "11"), -- i=1727
      ("1000011001100000", "00"), -- i=1728
      ("1001011001100000", "01"), -- i=1729
      ("1010011001100000", "10"), -- i=1730
      ("1011011001100000", "11"), -- i=1731
      ("1000011001100001", "00"), -- i=1732
      ("1001011001100001", "01"), -- i=1733
      ("1010011001100001", "10"), -- i=1734
      ("1011011001100001", "11"), -- i=1735
      ("1000011001100010", "00"), -- i=1736
      ("1001011001100010", "01"), -- i=1737
      ("1010011001100010", "10"), -- i=1738
      ("1011011001100010", "11"), -- i=1739
      ("1000011001100011", "00"), -- i=1740
      ("1001011001100011", "01"), -- i=1741
      ("1010011001100011", "10"), -- i=1742
      ("1011011001100011", "11"), -- i=1743
      ("1000011001100100", "00"), -- i=1744
      ("1001011001100100", "01"), -- i=1745
      ("1010011001100100", "10"), -- i=1746
      ("1011011001100100", "11"), -- i=1747
      ("1000011001100101", "00"), -- i=1748
      ("1001011001100101", "01"), -- i=1749
      ("1010011001100101", "10"), -- i=1750
      ("1011011001100101", "11"), -- i=1751
      ("1000011001100110", "00"), -- i=1752
      ("1001011001100110", "01"), -- i=1753
      ("1010011001100110", "10"), -- i=1754
      ("1011011001100110", "11"), -- i=1755
      ("1000011001100111", "00"), -- i=1756
      ("1001011001100111", "01"), -- i=1757
      ("1010011001100111", "10"), -- i=1758
      ("1011011001100111", "11"), -- i=1759
      ("1000011001110000", "00"), -- i=1760
      ("1001011001110000", "01"), -- i=1761
      ("1010011001110000", "10"), -- i=1762
      ("1011011001110000", "11"), -- i=1763
      ("1000011001110001", "00"), -- i=1764
      ("1001011001110001", "01"), -- i=1765
      ("1010011001110001", "10"), -- i=1766
      ("1011011001110001", "11"), -- i=1767
      ("1000011001110010", "00"), -- i=1768
      ("1001011001110010", "01"), -- i=1769
      ("1010011001110010", "10"), -- i=1770
      ("1011011001110010", "11"), -- i=1771
      ("1000011001110011", "00"), -- i=1772
      ("1001011001110011", "01"), -- i=1773
      ("1010011001110011", "10"), -- i=1774
      ("1011011001110011", "11"), -- i=1775
      ("1000011001110100", "00"), -- i=1776
      ("1001011001110100", "01"), -- i=1777
      ("1010011001110100", "10"), -- i=1778
      ("1011011001110100", "11"), -- i=1779
      ("1000011001110101", "00"), -- i=1780
      ("1001011001110101", "01"), -- i=1781
      ("1010011001110101", "10"), -- i=1782
      ("1011011001110101", "11"), -- i=1783
      ("1000011001110110", "00"), -- i=1784
      ("1001011001110110", "01"), -- i=1785
      ("1010011001110110", "10"), -- i=1786
      ("1011011001110110", "11"), -- i=1787
      ("1000011001110111", "00"), -- i=1788
      ("1001011001110111", "01"), -- i=1789
      ("1010011001110111", "10"), -- i=1790
      ("1011011001110111", "11"), -- i=1791
      ("1000011100000000", "00"), -- i=1792
      ("1001011100000000", "01"), -- i=1793
      ("1010011100000000", "10"), -- i=1794
      ("1011011100000000", "11"), -- i=1795
      ("1000011100000001", "00"), -- i=1796
      ("1001011100000001", "01"), -- i=1797
      ("1010011100000001", "10"), -- i=1798
      ("1011011100000001", "11"), -- i=1799
      ("1000011100000010", "00"), -- i=1800
      ("1001011100000010", "01"), -- i=1801
      ("1010011100000010", "10"), -- i=1802
      ("1011011100000010", "11"), -- i=1803
      ("1000011100000011", "00"), -- i=1804
      ("1001011100000011", "01"), -- i=1805
      ("1010011100000011", "10"), -- i=1806
      ("1011011100000011", "11"), -- i=1807
      ("1000011100000100", "00"), -- i=1808
      ("1001011100000100", "01"), -- i=1809
      ("1010011100000100", "10"), -- i=1810
      ("1011011100000100", "11"), -- i=1811
      ("1000011100000101", "00"), -- i=1812
      ("1001011100000101", "01"), -- i=1813
      ("1010011100000101", "10"), -- i=1814
      ("1011011100000101", "11"), -- i=1815
      ("1000011100000110", "00"), -- i=1816
      ("1001011100000110", "01"), -- i=1817
      ("1010011100000110", "10"), -- i=1818
      ("1011011100000110", "11"), -- i=1819
      ("1000011100000111", "00"), -- i=1820
      ("1001011100000111", "01"), -- i=1821
      ("1010011100000111", "10"), -- i=1822
      ("1011011100000111", "11"), -- i=1823
      ("1000011100010000", "00"), -- i=1824
      ("1001011100010000", "01"), -- i=1825
      ("1010011100010000", "10"), -- i=1826
      ("1011011100010000", "11"), -- i=1827
      ("1000011100010001", "00"), -- i=1828
      ("1001011100010001", "01"), -- i=1829
      ("1010011100010001", "10"), -- i=1830
      ("1011011100010001", "11"), -- i=1831
      ("1000011100010010", "00"), -- i=1832
      ("1001011100010010", "01"), -- i=1833
      ("1010011100010010", "10"), -- i=1834
      ("1011011100010010", "11"), -- i=1835
      ("1000011100010011", "00"), -- i=1836
      ("1001011100010011", "01"), -- i=1837
      ("1010011100010011", "10"), -- i=1838
      ("1011011100010011", "11"), -- i=1839
      ("1000011100010100", "00"), -- i=1840
      ("1001011100010100", "01"), -- i=1841
      ("1010011100010100", "10"), -- i=1842
      ("1011011100010100", "11"), -- i=1843
      ("1000011100010101", "00"), -- i=1844
      ("1001011100010101", "01"), -- i=1845
      ("1010011100010101", "10"), -- i=1846
      ("1011011100010101", "11"), -- i=1847
      ("1000011100010110", "00"), -- i=1848
      ("1001011100010110", "01"), -- i=1849
      ("1010011100010110", "10"), -- i=1850
      ("1011011100010110", "11"), -- i=1851
      ("1000011100010111", "00"), -- i=1852
      ("1001011100010111", "01"), -- i=1853
      ("1010011100010111", "10"), -- i=1854
      ("1011011100010111", "11"), -- i=1855
      ("1000011100100000", "00"), -- i=1856
      ("1001011100100000", "01"), -- i=1857
      ("1010011100100000", "10"), -- i=1858
      ("1011011100100000", "11"), -- i=1859
      ("1000011100100001", "00"), -- i=1860
      ("1001011100100001", "01"), -- i=1861
      ("1010011100100001", "10"), -- i=1862
      ("1011011100100001", "11"), -- i=1863
      ("1000011100100010", "00"), -- i=1864
      ("1001011100100010", "01"), -- i=1865
      ("1010011100100010", "10"), -- i=1866
      ("1011011100100010", "11"), -- i=1867
      ("1000011100100011", "00"), -- i=1868
      ("1001011100100011", "01"), -- i=1869
      ("1010011100100011", "10"), -- i=1870
      ("1011011100100011", "11"), -- i=1871
      ("1000011100100100", "00"), -- i=1872
      ("1001011100100100", "01"), -- i=1873
      ("1010011100100100", "10"), -- i=1874
      ("1011011100100100", "11"), -- i=1875
      ("1000011100100101", "00"), -- i=1876
      ("1001011100100101", "01"), -- i=1877
      ("1010011100100101", "10"), -- i=1878
      ("1011011100100101", "11"), -- i=1879
      ("1000011100100110", "00"), -- i=1880
      ("1001011100100110", "01"), -- i=1881
      ("1010011100100110", "10"), -- i=1882
      ("1011011100100110", "11"), -- i=1883
      ("1000011100100111", "00"), -- i=1884
      ("1001011100100111", "01"), -- i=1885
      ("1010011100100111", "10"), -- i=1886
      ("1011011100100111", "11"), -- i=1887
      ("1000011100110000", "00"), -- i=1888
      ("1001011100110000", "01"), -- i=1889
      ("1010011100110000", "10"), -- i=1890
      ("1011011100110000", "11"), -- i=1891
      ("1000011100110001", "00"), -- i=1892
      ("1001011100110001", "01"), -- i=1893
      ("1010011100110001", "10"), -- i=1894
      ("1011011100110001", "11"), -- i=1895
      ("1000011100110010", "00"), -- i=1896
      ("1001011100110010", "01"), -- i=1897
      ("1010011100110010", "10"), -- i=1898
      ("1011011100110010", "11"), -- i=1899
      ("1000011100110011", "00"), -- i=1900
      ("1001011100110011", "01"), -- i=1901
      ("1010011100110011", "10"), -- i=1902
      ("1011011100110011", "11"), -- i=1903
      ("1000011100110100", "00"), -- i=1904
      ("1001011100110100", "01"), -- i=1905
      ("1010011100110100", "10"), -- i=1906
      ("1011011100110100", "11"), -- i=1907
      ("1000011100110101", "00"), -- i=1908
      ("1001011100110101", "01"), -- i=1909
      ("1010011100110101", "10"), -- i=1910
      ("1011011100110101", "11"), -- i=1911
      ("1000011100110110", "00"), -- i=1912
      ("1001011100110110", "01"), -- i=1913
      ("1010011100110110", "10"), -- i=1914
      ("1011011100110110", "11"), -- i=1915
      ("1000011100110111", "00"), -- i=1916
      ("1001011100110111", "01"), -- i=1917
      ("1010011100110111", "10"), -- i=1918
      ("1011011100110111", "11"), -- i=1919
      ("1000011101000000", "00"), -- i=1920
      ("1001011101000000", "01"), -- i=1921
      ("1010011101000000", "10"), -- i=1922
      ("1011011101000000", "11"), -- i=1923
      ("1000011101000001", "00"), -- i=1924
      ("1001011101000001", "01"), -- i=1925
      ("1010011101000001", "10"), -- i=1926
      ("1011011101000001", "11"), -- i=1927
      ("1000011101000010", "00"), -- i=1928
      ("1001011101000010", "01"), -- i=1929
      ("1010011101000010", "10"), -- i=1930
      ("1011011101000010", "11"), -- i=1931
      ("1000011101000011", "00"), -- i=1932
      ("1001011101000011", "01"), -- i=1933
      ("1010011101000011", "10"), -- i=1934
      ("1011011101000011", "11"), -- i=1935
      ("1000011101000100", "00"), -- i=1936
      ("1001011101000100", "01"), -- i=1937
      ("1010011101000100", "10"), -- i=1938
      ("1011011101000100", "11"), -- i=1939
      ("1000011101000101", "00"), -- i=1940
      ("1001011101000101", "01"), -- i=1941
      ("1010011101000101", "10"), -- i=1942
      ("1011011101000101", "11"), -- i=1943
      ("1000011101000110", "00"), -- i=1944
      ("1001011101000110", "01"), -- i=1945
      ("1010011101000110", "10"), -- i=1946
      ("1011011101000110", "11"), -- i=1947
      ("1000011101000111", "00"), -- i=1948
      ("1001011101000111", "01"), -- i=1949
      ("1010011101000111", "10"), -- i=1950
      ("1011011101000111", "11"), -- i=1951
      ("1000011101010000", "00"), -- i=1952
      ("1001011101010000", "01"), -- i=1953
      ("1010011101010000", "10"), -- i=1954
      ("1011011101010000", "11"), -- i=1955
      ("1000011101010001", "00"), -- i=1956
      ("1001011101010001", "01"), -- i=1957
      ("1010011101010001", "10"), -- i=1958
      ("1011011101010001", "11"), -- i=1959
      ("1000011101010010", "00"), -- i=1960
      ("1001011101010010", "01"), -- i=1961
      ("1010011101010010", "10"), -- i=1962
      ("1011011101010010", "11"), -- i=1963
      ("1000011101010011", "00"), -- i=1964
      ("1001011101010011", "01"), -- i=1965
      ("1010011101010011", "10"), -- i=1966
      ("1011011101010011", "11"), -- i=1967
      ("1000011101010100", "00"), -- i=1968
      ("1001011101010100", "01"), -- i=1969
      ("1010011101010100", "10"), -- i=1970
      ("1011011101010100", "11"), -- i=1971
      ("1000011101010101", "00"), -- i=1972
      ("1001011101010101", "01"), -- i=1973
      ("1010011101010101", "10"), -- i=1974
      ("1011011101010101", "11"), -- i=1975
      ("1000011101010110", "00"), -- i=1976
      ("1001011101010110", "01"), -- i=1977
      ("1010011101010110", "10"), -- i=1978
      ("1011011101010110", "11"), -- i=1979
      ("1000011101010111", "00"), -- i=1980
      ("1001011101010111", "01"), -- i=1981
      ("1010011101010111", "10"), -- i=1982
      ("1011011101010111", "11"), -- i=1983
      ("1000011101100000", "00"), -- i=1984
      ("1001011101100000", "01"), -- i=1985
      ("1010011101100000", "10"), -- i=1986
      ("1011011101100000", "11"), -- i=1987
      ("1000011101100001", "00"), -- i=1988
      ("1001011101100001", "01"), -- i=1989
      ("1010011101100001", "10"), -- i=1990
      ("1011011101100001", "11"), -- i=1991
      ("1000011101100010", "00"), -- i=1992
      ("1001011101100010", "01"), -- i=1993
      ("1010011101100010", "10"), -- i=1994
      ("1011011101100010", "11"), -- i=1995
      ("1000011101100011", "00"), -- i=1996
      ("1001011101100011", "01"), -- i=1997
      ("1010011101100011", "10"), -- i=1998
      ("1011011101100011", "11"), -- i=1999
      ("1000011101100100", "00"), -- i=2000
      ("1001011101100100", "01"), -- i=2001
      ("1010011101100100", "10"), -- i=2002
      ("1011011101100100", "11"), -- i=2003
      ("1000011101100101", "00"), -- i=2004
      ("1001011101100101", "01"), -- i=2005
      ("1010011101100101", "10"), -- i=2006
      ("1011011101100101", "11"), -- i=2007
      ("1000011101100110", "00"), -- i=2008
      ("1001011101100110", "01"), -- i=2009
      ("1010011101100110", "10"), -- i=2010
      ("1011011101100110", "11"), -- i=2011
      ("1000011101100111", "00"), -- i=2012
      ("1001011101100111", "01"), -- i=2013
      ("1010011101100111", "10"), -- i=2014
      ("1011011101100111", "11"), -- i=2015
      ("1000011101110000", "00"), -- i=2016
      ("1001011101110000", "01"), -- i=2017
      ("1010011101110000", "10"), -- i=2018
      ("1011011101110000", "11"), -- i=2019
      ("1000011101110001", "00"), -- i=2020
      ("1001011101110001", "01"), -- i=2021
      ("1010011101110001", "10"), -- i=2022
      ("1011011101110001", "11"), -- i=2023
      ("1000011101110010", "00"), -- i=2024
      ("1001011101110010", "01"), -- i=2025
      ("1010011101110010", "10"), -- i=2026
      ("1011011101110010", "11"), -- i=2027
      ("1000011101110011", "00"), -- i=2028
      ("1001011101110011", "01"), -- i=2029
      ("1010011101110011", "10"), -- i=2030
      ("1011011101110011", "11"), -- i=2031
      ("1000011101110100", "00"), -- i=2032
      ("1001011101110100", "01"), -- i=2033
      ("1010011101110100", "10"), -- i=2034
      ("1011011101110100", "11"), -- i=2035
      ("1000011101110101", "00"), -- i=2036
      ("1001011101110101", "01"), -- i=2037
      ("1010011101110101", "10"), -- i=2038
      ("1011011101110101", "11"), -- i=2039
      ("1000011101110110", "00"), -- i=2040
      ("1001011101110110", "01"), -- i=2041
      ("1010011101110110", "10"), -- i=2042
      ("1011011101110110", "11"), -- i=2043
      ("1000011101110111", "00"), -- i=2044
      ("1001011101110111", "01"), -- i=2045
      ("1010011101110111", "10"), -- i=2046
      ("1011011101110111", "11"));
  begin
    for i in patterns'range loop
      INST <= patterns(i).INST;
      FL_Z <= patterns(i).FL_Z;
      wait for 10 ns;
      assert std_match(ALUOP, patterns(i).ALUOP) OR (ALUOP = "ZZ" AND patterns(i).ALUOP = "ZZ")
        report "wrong value for ALUOP, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).ALUOP) & ", found " & to_string(ALUOP) severity error;assert std_match(RS1, patterns(i).RS1) OR (RS1 = "ZZZ" AND patterns(i).RS1 = "ZZZ")
        report "wrong value for RS1, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).RS1) & ", found " & to_string(RS1) severity error;assert std_match(RS2, patterns(i).RS2) OR (RS2 = "ZZZ" AND patterns(i).RS2 = "ZZZ")
        report "wrong value for RS2, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).RS2) & ", found " & to_string(RS2) severity error;assert std_match(WS, patterns(i).WS) OR (WS = "ZZZ" AND patterns(i).WS = "ZZZ")
        report "wrong value for WS, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).WS) & ", found " & to_string(WS) severity error;assert std_match(STR, patterns(i).STR) OR (STR = 'Z' AND patterns(i).STR = 'Z')
        report "wrong value for STR, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).STR) & ", found " & std_logic'image(STR) severity error;assert std_match(WE, patterns(i).WE) OR (WE = 'Z' AND patterns(i).WE = 'Z')
        report "wrong value for WE, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).WE) & ", found " & std_logic'image(WE) severity error;assert std_match(DMUX, patterns(i).DMUX) OR (DMUX = "ZZ" AND patterns(i).DMUX = "ZZ")
        report "wrong value for DMUX, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).DMUX) & ", found " & to_string(DMUX) severity error;assert std_match(LDR, patterns(i).LDR) OR (LDR = 'Z' AND patterns(i).LDR = 'Z')
        report "wrong value for LDR, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).LDR) & ", found " & std_logic'image(LDR) severity error;assert std_match(FL_EN, patterns(i).FL_EN) OR (FL_EN = 'Z' AND patterns(i).FL_EN = 'Z')
        report "wrong value for FL_EN, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).FL_EN) & ", found " & std_logic'image(FL_EN) severity error;assert std_match(HE, patterns(i).HE) OR (HE = 'Z' AND patterns(i).HE = 'Z')
        report "wrong value for HE, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).HE) & ", found " & std_logic'image(HE) severity error;end loop;
    wait;
  end process;
end behav;
