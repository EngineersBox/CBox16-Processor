--  A testbench for control_unit_All_Tests_tb
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity control_unit_All_Tests_tb is
end control_unit_All_Tests_tb;

architecture behav of control_unit_All_Tests_tb is
  component main
    port (
      INST: in std_logic_vector(15 downto 0);
      FL_Z: in std_logic;
      ALUOP: out std_logic_vector(1 downto 0);
      RS1: out std_logic_vector(2 downto 0);
      RS2: out std_logic_vector(2 downto 0);
      WS: out std_logic_vector(2 downto 0);
      STR: out std_logic;
      WE: out std_logic;
      DMUX: out std_logic_vector(1 downto 0);
      LDR: out std_logic;
      FL_EN: out std_logic;
      HE: out std_logic);
  end component;

  signal INST : std_logic_vector(15 downto 0);
  signal FL_Z : std_logic;
  signal ALUOP : std_logic_vector(1 downto 0);
  signal RS1 : std_logic_vector(2 downto 0);
  signal RS2 : std_logic_vector(2 downto 0);
  signal WS : std_logic_vector(2 downto 0);
  signal STR : std_logic;
  signal WE : std_logic;
  signal DMUX : std_logic_vector(1 downto 0);
  signal LDR : std_logic;
  signal FL_EN : std_logic;
  signal HE : std_logic;
  function to_string ( a: std_logic_vector) return string is
      variable b : string (1 to a'length) := (others => NUL);
      variable stri : integer := 1; 
  begin
      for i in a'range loop
          b(stri) := std_logic'image(a((i)))(2);
      stri := stri+1;
      end loop;
      return b;
  end function;
begin
  main_0 : main port map (
    INST => INST,
    FL_Z => FL_Z,
    ALUOP => ALUOP,
    RS1 => RS1,
    RS2 => RS2,
    WS => WS,
    STR => STR,
    WE => WE,
    DMUX => DMUX,
    LDR => LDR,
    FL_EN => FL_EN,
    HE => HE );
  process
    type pattern_type is record
      INST : std_logic_vector(15 downto 0);
      FL_Z : std_logic;
      WE : std_logic;
      ALUOP : std_logic_vector(1 downto 0);
      RS1 : std_logic_vector(2 downto 0);
      RS2 : std_logic_vector(2 downto 0);
      WS : std_logic_vector(2 downto 0);
      STR : std_logic;
      LDR : std_logic;
      DMUX : std_logic_vector(1 downto 0);
    end record;
    type pattern_array is array (natural range <>) of pattern_type;
    constant patterns : pattern_array := (
      ("1000000000000000", '0', '1', "00", "000", "000", "000", '0', '-', "00"), -- i=0
      ("1000100000000000", '1', '1', "00", "000", "000", "000", '0', '-', "00"), -- i=1
      ("1000100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2
      ("1001000000000000", '0', '1', "01", "000", "000", "000", '0', '-', "00"), -- i=3
      ("1001100000000000", '1', '1', "01", "000", "000", "000", '0', '-', "00"), -- i=4
      ("1001100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5
      ("1010000000000000", '0', '1', "10", "000", "000", "000", '0', '-', "00"), -- i=6
      ("1010100000000000", '1', '1', "10", "000", "000", "000", '0', '-', "00"), -- i=7
      ("1010100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8
      ("1011000000000000", '0', '1', "11", "000", "000", "000", '0', '-', "00"), -- i=9
      ("1011100000000000", '1', '1', "11", "000", "000", "000", '0', '-', "00"), -- i=10
      ("1011100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=11
      ("0101000000000000", '0', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=12
      ("0101100000000000", '1', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=13
      ("0101100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=14
      ("0100000000000000", '0', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=15
      ("0100100000000000", '1', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=16
      ("0100100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=17
      ("0000000000001101", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=18
      ("0000100000001101", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=19
      ("0000100000001101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=20
      ("1000000000000001", '0', '1', "00", "000", "001", "000", '0', '-', "00"), -- i=21
      ("1000100000000001", '1', '1', "00", "000", "001", "000", '0', '-', "00"), -- i=22
      ("1000100000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=23
      ("1001000000000001", '0', '1', "01", "000", "001", "000", '0', '-', "00"), -- i=24
      ("1001100000000001", '1', '1', "01", "000", "001", "000", '0', '-', "00"), -- i=25
      ("1001100000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=26
      ("1010000000000001", '0', '1', "10", "000", "001", "000", '0', '-', "00"), -- i=27
      ("1010100000000001", '1', '1', "10", "000", "001", "000", '0', '-', "00"), -- i=28
      ("1010100000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=29
      ("1011000000000001", '0', '1', "11", "000", "001", "000", '0', '-', "00"), -- i=30
      ("1011100000000001", '1', '1', "11", "000", "001", "000", '0', '-', "00"), -- i=31
      ("1011100000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=32
      ("0101000000000000", '0', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=33
      ("0101100000000000", '1', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=34
      ("0101100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=35
      ("0100000000000000", '0', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=36
      ("0100100000000000", '1', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=37
      ("0100100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=38
      ("0000000010010101", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=39
      ("0000100010010101", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=40
      ("0000100010010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=41
      ("1000000000000010", '0', '1', "00", "000", "010", "000", '0', '-', "00"), -- i=42
      ("1000100000000010", '1', '1', "00", "000", "010", "000", '0', '-', "00"), -- i=43
      ("1000100000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=44
      ("1001000000000010", '0', '1', "01", "000", "010", "000", '0', '-', "00"), -- i=45
      ("1001100000000010", '1', '1', "01", "000", "010", "000", '0', '-', "00"), -- i=46
      ("1001100000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=47
      ("1010000000000010", '0', '1', "10", "000", "010", "000", '0', '-', "00"), -- i=48
      ("1010100000000010", '1', '1', "10", "000", "010", "000", '0', '-', "00"), -- i=49
      ("1010100000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=50
      ("1011000000000010", '0', '1', "11", "000", "010", "000", '0', '-', "00"), -- i=51
      ("1011100000000010", '1', '1', "11", "000", "010", "000", '0', '-', "00"), -- i=52
      ("1011100000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=53
      ("0101000000000000", '0', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=54
      ("0101100000000000", '1', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=55
      ("0101100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=56
      ("0100000000000000", '0', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=57
      ("0100100000000000", '1', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=58
      ("0100100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=59
      ("0000000001000010", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=60
      ("0000100001000010", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=61
      ("0000100001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=62
      ("1000000000000011", '0', '1', "00", "000", "011", "000", '0', '-', "00"), -- i=63
      ("1000100000000011", '1', '1', "00", "000", "011", "000", '0', '-', "00"), -- i=64
      ("1000100000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=65
      ("1001000000000011", '0', '1', "01", "000", "011", "000", '0', '-', "00"), -- i=66
      ("1001100000000011", '1', '1', "01", "000", "011", "000", '0', '-', "00"), -- i=67
      ("1001100000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=68
      ("1010000000000011", '0', '1', "10", "000", "011", "000", '0', '-', "00"), -- i=69
      ("1010100000000011", '1', '1', "10", "000", "011", "000", '0', '-', "00"), -- i=70
      ("1010100000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=71
      ("1011000000000011", '0', '1', "11", "000", "011", "000", '0', '-', "00"), -- i=72
      ("1011100000000011", '1', '1', "11", "000", "011", "000", '0', '-', "00"), -- i=73
      ("1011100000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=74
      ("0101000000000000", '0', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=75
      ("0101100000000000", '1', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=76
      ("0101100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=77
      ("0100000000000000", '0', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=78
      ("0100100000000000", '1', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=79
      ("0100100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=80
      ("0000000010110001", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=81
      ("0000100010110001", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=82
      ("0000100010110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=83
      ("1000000000000100", '0', '1', "00", "000", "100", "000", '0', '-', "00"), -- i=84
      ("1000100000000100", '1', '1', "00", "000", "100", "000", '0', '-', "00"), -- i=85
      ("1000100000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=86
      ("1001000000000100", '0', '1', "01", "000", "100", "000", '0', '-', "00"), -- i=87
      ("1001100000000100", '1', '1', "01", "000", "100", "000", '0', '-', "00"), -- i=88
      ("1001100000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=89
      ("1010000000000100", '0', '1', "10", "000", "100", "000", '0', '-', "00"), -- i=90
      ("1010100000000100", '1', '1', "10", "000", "100", "000", '0', '-', "00"), -- i=91
      ("1010100000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=92
      ("1011000000000100", '0', '1', "11", "000", "100", "000", '0', '-', "00"), -- i=93
      ("1011100000000100", '1', '1', "11", "000", "100", "000", '0', '-', "00"), -- i=94
      ("1011100000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=95
      ("0101000000000000", '0', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=96
      ("0101100000000000", '1', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=97
      ("0101100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=98
      ("0100000000000000", '0', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=99
      ("0100100000000000", '1', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=100
      ("0100100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=101
      ("0000000001110100", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=102
      ("0000100001110100", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=103
      ("0000100001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=104
      ("1000000000000101", '0', '1', "00", "000", "101", "000", '0', '-', "00"), -- i=105
      ("1000100000000101", '1', '1', "00", "000", "101", "000", '0', '-', "00"), -- i=106
      ("1000100000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=107
      ("1001000000000101", '0', '1', "01", "000", "101", "000", '0', '-', "00"), -- i=108
      ("1001100000000101", '1', '1', "01", "000", "101", "000", '0', '-', "00"), -- i=109
      ("1001100000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=110
      ("1010000000000101", '0', '1', "10", "000", "101", "000", '0', '-', "00"), -- i=111
      ("1010100000000101", '1', '1', "10", "000", "101", "000", '0', '-', "00"), -- i=112
      ("1010100000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=113
      ("1011000000000101", '0', '1', "11", "000", "101", "000", '0', '-', "00"), -- i=114
      ("1011100000000101", '1', '1', "11", "000", "101", "000", '0', '-', "00"), -- i=115
      ("1011100000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=116
      ("0101000000000000", '0', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=117
      ("0101100000000000", '1', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=118
      ("0101100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=119
      ("0100000000000000", '0', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=120
      ("0100100000000000", '1', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=121
      ("0100100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=122
      ("0000000011001101", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=123
      ("0000100011001101", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=124
      ("0000100011001101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=125
      ("1000000000000110", '0', '1', "00", "000", "110", "000", '0', '-', "00"), -- i=126
      ("1000100000000110", '1', '1', "00", "000", "110", "000", '0', '-', "00"), -- i=127
      ("1000100000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=128
      ("1001000000000110", '0', '1', "01", "000", "110", "000", '0', '-', "00"), -- i=129
      ("1001100000000110", '1', '1', "01", "000", "110", "000", '0', '-', "00"), -- i=130
      ("1001100000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=131
      ("1010000000000110", '0', '1', "10", "000", "110", "000", '0', '-', "00"), -- i=132
      ("1010100000000110", '1', '1', "10", "000", "110", "000", '0', '-', "00"), -- i=133
      ("1010100000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=134
      ("1011000000000110", '0', '1', "11", "000", "110", "000", '0', '-', "00"), -- i=135
      ("1011100000000110", '1', '1', "11", "000", "110", "000", '0', '-', "00"), -- i=136
      ("1011100000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=137
      ("0101000000000000", '0', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=138
      ("0101100000000000", '1', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=139
      ("0101100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=140
      ("0100000000000000", '0', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=141
      ("0100100000000000", '1', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=142
      ("0100100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=143
      ("0000000000110100", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=144
      ("0000100000110100", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=145
      ("0000100000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=146
      ("1000000000000111", '0', '1', "00", "000", "111", "000", '0', '-', "00"), -- i=147
      ("1000100000000111", '1', '1', "00", "000", "111", "000", '0', '-', "00"), -- i=148
      ("1000100000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=149
      ("1001000000000111", '0', '1', "01", "000", "111", "000", '0', '-', "00"), -- i=150
      ("1001100000000111", '1', '1', "01", "000", "111", "000", '0', '-', "00"), -- i=151
      ("1001100000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=152
      ("1010000000000111", '0', '1', "10", "000", "111", "000", '0', '-', "00"), -- i=153
      ("1010100000000111", '1', '1', "10", "000", "111", "000", '0', '-', "00"), -- i=154
      ("1010100000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=155
      ("1011000000000111", '0', '1', "11", "000", "111", "000", '0', '-', "00"), -- i=156
      ("1011100000000111", '1', '1', "11", "000", "111", "000", '0', '-', "00"), -- i=157
      ("1011100000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=158
      ("0101000000000000", '0', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=159
      ("0101100000000000", '1', '1', "--", "000", "---", "000", '0', '1', "01"), -- i=160
      ("0101100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=161
      ("0100000000000000", '0', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=162
      ("0100100000000000", '1', '0', "--", "000", "000", "---", '1', '-', "--"), -- i=163
      ("0100100000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=164
      ("0000000010110111", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=165
      ("0000100010110111", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=166
      ("0000100010110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=167
      ("1000000000010000", '0', '1', "00", "001", "000", "000", '0', '-', "00"), -- i=168
      ("1000100000010000", '1', '1', "00", "001", "000", "000", '0', '-', "00"), -- i=169
      ("1000100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=170
      ("1001000000010000", '0', '1', "01", "001", "000", "000", '0', '-', "00"), -- i=171
      ("1001100000010000", '1', '1', "01", "001", "000", "000", '0', '-', "00"), -- i=172
      ("1001100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=173
      ("1010000000010000", '0', '1', "10", "001", "000", "000", '0', '-', "00"), -- i=174
      ("1010100000010000", '1', '1', "10", "001", "000", "000", '0', '-', "00"), -- i=175
      ("1010100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=176
      ("1011000000010000", '0', '1', "11", "001", "000", "000", '0', '-', "00"), -- i=177
      ("1011100000010000", '1', '1', "11", "001", "000", "000", '0', '-', "00"), -- i=178
      ("1011100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=179
      ("0101000000010000", '0', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=180
      ("0101100000010000", '1', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=181
      ("0101100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=182
      ("0100000000010000", '0', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=183
      ("0100100000010000", '1', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=184
      ("0100100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=185
      ("0000000010011010", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=186
      ("0000100010011010", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=187
      ("0000100010011010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=188
      ("1000000000010001", '0', '1', "00", "001", "001", "000", '0', '-', "00"), -- i=189
      ("1000100000010001", '1', '1', "00", "001", "001", "000", '0', '-', "00"), -- i=190
      ("1000100000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=191
      ("1001000000010001", '0', '1', "01", "001", "001", "000", '0', '-', "00"), -- i=192
      ("1001100000010001", '1', '1', "01", "001", "001", "000", '0', '-', "00"), -- i=193
      ("1001100000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=194
      ("1010000000010001", '0', '1', "10", "001", "001", "000", '0', '-', "00"), -- i=195
      ("1010100000010001", '1', '1', "10", "001", "001", "000", '0', '-', "00"), -- i=196
      ("1010100000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=197
      ("1011000000010001", '0', '1', "11", "001", "001", "000", '0', '-', "00"), -- i=198
      ("1011100000010001", '1', '1', "11", "001", "001", "000", '0', '-', "00"), -- i=199
      ("1011100000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=200
      ("0101000000010000", '0', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=201
      ("0101100000010000", '1', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=202
      ("0101100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=203
      ("0100000000010000", '0', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=204
      ("0100100000010000", '1', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=205
      ("0100100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=206
      ("0000000011110111", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=207
      ("0000100011110111", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=208
      ("0000100011110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=209
      ("1000000000010010", '0', '1', "00", "001", "010", "000", '0', '-', "00"), -- i=210
      ("1000100000010010", '1', '1', "00", "001", "010", "000", '0', '-', "00"), -- i=211
      ("1000100000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=212
      ("1001000000010010", '0', '1', "01", "001", "010", "000", '0', '-', "00"), -- i=213
      ("1001100000010010", '1', '1', "01", "001", "010", "000", '0', '-', "00"), -- i=214
      ("1001100000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=215
      ("1010000000010010", '0', '1', "10", "001", "010", "000", '0', '-', "00"), -- i=216
      ("1010100000010010", '1', '1', "10", "001", "010", "000", '0', '-', "00"), -- i=217
      ("1010100000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=218
      ("1011000000010010", '0', '1', "11", "001", "010", "000", '0', '-', "00"), -- i=219
      ("1011100000010010", '1', '1', "11", "001", "010", "000", '0', '-', "00"), -- i=220
      ("1011100000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=221
      ("0101000000010000", '0', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=222
      ("0101100000010000", '1', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=223
      ("0101100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=224
      ("0100000000010000", '0', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=225
      ("0100100000010000", '1', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=226
      ("0100100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=227
      ("0000000001001101", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=228
      ("0000100001001101", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=229
      ("0000100001001101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=230
      ("1000000000010011", '0', '1', "00", "001", "011", "000", '0', '-', "00"), -- i=231
      ("1000100000010011", '1', '1', "00", "001", "011", "000", '0', '-', "00"), -- i=232
      ("1000100000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=233
      ("1001000000010011", '0', '1', "01", "001", "011", "000", '0', '-', "00"), -- i=234
      ("1001100000010011", '1', '1', "01", "001", "011", "000", '0', '-', "00"), -- i=235
      ("1001100000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=236
      ("1010000000010011", '0', '1', "10", "001", "011", "000", '0', '-', "00"), -- i=237
      ("1010100000010011", '1', '1', "10", "001", "011", "000", '0', '-', "00"), -- i=238
      ("1010100000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=239
      ("1011000000010011", '0', '1', "11", "001", "011", "000", '0', '-', "00"), -- i=240
      ("1011100000010011", '1', '1', "11", "001", "011", "000", '0', '-', "00"), -- i=241
      ("1011100000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=242
      ("0101000000010000", '0', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=243
      ("0101100000010000", '1', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=244
      ("0101100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=245
      ("0100000000010000", '0', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=246
      ("0100100000010000", '1', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=247
      ("0100100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=248
      ("0000000001000010", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=249
      ("0000100001000010", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=250
      ("0000100001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=251
      ("1000000000010100", '0', '1', "00", "001", "100", "000", '0', '-', "00"), -- i=252
      ("1000100000010100", '1', '1', "00", "001", "100", "000", '0', '-', "00"), -- i=253
      ("1000100000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=254
      ("1001000000010100", '0', '1', "01", "001", "100", "000", '0', '-', "00"), -- i=255
      ("1001100000010100", '1', '1', "01", "001", "100", "000", '0', '-', "00"), -- i=256
      ("1001100000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=257
      ("1010000000010100", '0', '1', "10", "001", "100", "000", '0', '-', "00"), -- i=258
      ("1010100000010100", '1', '1', "10", "001", "100", "000", '0', '-', "00"), -- i=259
      ("1010100000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=260
      ("1011000000010100", '0', '1', "11", "001", "100", "000", '0', '-', "00"), -- i=261
      ("1011100000010100", '1', '1', "11", "001", "100", "000", '0', '-', "00"), -- i=262
      ("1011100000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=263
      ("0101000000010000", '0', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=264
      ("0101100000010000", '1', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=265
      ("0101100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=266
      ("0100000000010000", '0', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=267
      ("0100100000010000", '1', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=268
      ("0100100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=269
      ("0000000010010111", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=270
      ("0000100010010111", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=271
      ("0000100010010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=272
      ("1000000000010101", '0', '1', "00", "001", "101", "000", '0', '-', "00"), -- i=273
      ("1000100000010101", '1', '1', "00", "001", "101", "000", '0', '-', "00"), -- i=274
      ("1000100000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=275
      ("1001000000010101", '0', '1', "01", "001", "101", "000", '0', '-', "00"), -- i=276
      ("1001100000010101", '1', '1', "01", "001", "101", "000", '0', '-', "00"), -- i=277
      ("1001100000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=278
      ("1010000000010101", '0', '1', "10", "001", "101", "000", '0', '-', "00"), -- i=279
      ("1010100000010101", '1', '1', "10", "001", "101", "000", '0', '-', "00"), -- i=280
      ("1010100000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=281
      ("1011000000010101", '0', '1', "11", "001", "101", "000", '0', '-', "00"), -- i=282
      ("1011100000010101", '1', '1', "11", "001", "101", "000", '0', '-', "00"), -- i=283
      ("1011100000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=284
      ("0101000000010000", '0', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=285
      ("0101100000010000", '1', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=286
      ("0101100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=287
      ("0100000000010000", '0', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=288
      ("0100100000010000", '1', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=289
      ("0100100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=290
      ("0000000011001100", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=291
      ("0000100011001100", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=292
      ("0000100011001100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=293
      ("1000000000010110", '0', '1', "00", "001", "110", "000", '0', '-', "00"), -- i=294
      ("1000100000010110", '1', '1', "00", "001", "110", "000", '0', '-', "00"), -- i=295
      ("1000100000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=296
      ("1001000000010110", '0', '1', "01", "001", "110", "000", '0', '-', "00"), -- i=297
      ("1001100000010110", '1', '1', "01", "001", "110", "000", '0', '-', "00"), -- i=298
      ("1001100000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=299
      ("1010000000010110", '0', '1', "10", "001", "110", "000", '0', '-', "00"), -- i=300
      ("1010100000010110", '1', '1', "10", "001", "110", "000", '0', '-', "00"), -- i=301
      ("1010100000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=302
      ("1011000000010110", '0', '1', "11", "001", "110", "000", '0', '-', "00"), -- i=303
      ("1011100000010110", '1', '1', "11", "001", "110", "000", '0', '-', "00"), -- i=304
      ("1011100000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=305
      ("0101000000010000", '0', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=306
      ("0101100000010000", '1', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=307
      ("0101100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=308
      ("0100000000010000", '0', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=309
      ("0100100000010000", '1', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=310
      ("0100100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=311
      ("0000000000100100", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=312
      ("0000100000100100", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=313
      ("0000100000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=314
      ("1000000000010111", '0', '1', "00", "001", "111", "000", '0', '-', "00"), -- i=315
      ("1000100000010111", '1', '1', "00", "001", "111", "000", '0', '-', "00"), -- i=316
      ("1000100000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=317
      ("1001000000010111", '0', '1', "01", "001", "111", "000", '0', '-', "00"), -- i=318
      ("1001100000010111", '1', '1', "01", "001", "111", "000", '0', '-', "00"), -- i=319
      ("1001100000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=320
      ("1010000000010111", '0', '1', "10", "001", "111", "000", '0', '-', "00"), -- i=321
      ("1010100000010111", '1', '1', "10", "001", "111", "000", '0', '-', "00"), -- i=322
      ("1010100000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=323
      ("1011000000010111", '0', '1', "11", "001", "111", "000", '0', '-', "00"), -- i=324
      ("1011100000010111", '1', '1', "11", "001", "111", "000", '0', '-', "00"), -- i=325
      ("1011100000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=326
      ("0101000000010000", '0', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=327
      ("0101100000010000", '1', '1', "--", "001", "---", "000", '0', '1', "01"), -- i=328
      ("0101100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=329
      ("0100000000010000", '0', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=330
      ("0100100000010000", '1', '0', "--", "001", "000", "---", '1', '-', "--"), -- i=331
      ("0100100000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=332
      ("0000000001100101", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=333
      ("0000100001100101", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=334
      ("0000100001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=335
      ("1000000000100000", '0', '1', "00", "010", "000", "000", '0', '-', "00"), -- i=336
      ("1000100000100000", '1', '1', "00", "010", "000", "000", '0', '-', "00"), -- i=337
      ("1000100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=338
      ("1001000000100000", '0', '1', "01", "010", "000", "000", '0', '-', "00"), -- i=339
      ("1001100000100000", '1', '1', "01", "010", "000", "000", '0', '-', "00"), -- i=340
      ("1001100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=341
      ("1010000000100000", '0', '1', "10", "010", "000", "000", '0', '-', "00"), -- i=342
      ("1010100000100000", '1', '1', "10", "010", "000", "000", '0', '-', "00"), -- i=343
      ("1010100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=344
      ("1011000000100000", '0', '1', "11", "010", "000", "000", '0', '-', "00"), -- i=345
      ("1011100000100000", '1', '1', "11", "010", "000", "000", '0', '-', "00"), -- i=346
      ("1011100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=347
      ("0101000000100000", '0', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=348
      ("0101100000100000", '1', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=349
      ("0101100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=350
      ("0100000000100000", '0', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=351
      ("0100100000100000", '1', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=352
      ("0100100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=353
      ("0000000011110001", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=354
      ("0000100011110001", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=355
      ("0000100011110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=356
      ("1000000000100001", '0', '1', "00", "010", "001", "000", '0', '-', "00"), -- i=357
      ("1000100000100001", '1', '1', "00", "010", "001", "000", '0', '-', "00"), -- i=358
      ("1000100000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=359
      ("1001000000100001", '0', '1', "01", "010", "001", "000", '0', '-', "00"), -- i=360
      ("1001100000100001", '1', '1', "01", "010", "001", "000", '0', '-', "00"), -- i=361
      ("1001100000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=362
      ("1010000000100001", '0', '1', "10", "010", "001", "000", '0', '-', "00"), -- i=363
      ("1010100000100001", '1', '1', "10", "010", "001", "000", '0', '-', "00"), -- i=364
      ("1010100000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=365
      ("1011000000100001", '0', '1', "11", "010", "001", "000", '0', '-', "00"), -- i=366
      ("1011100000100001", '1', '1', "11", "010", "001", "000", '0', '-', "00"), -- i=367
      ("1011100000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=368
      ("0101000000100000", '0', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=369
      ("0101100000100000", '1', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=370
      ("0101100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=371
      ("0100000000100000", '0', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=372
      ("0100100000100000", '1', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=373
      ("0100100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=374
      ("0000000001010110", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=375
      ("0000100001010110", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=376
      ("0000100001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=377
      ("1000000000100010", '0', '1', "00", "010", "010", "000", '0', '-', "00"), -- i=378
      ("1000100000100010", '1', '1', "00", "010", "010", "000", '0', '-', "00"), -- i=379
      ("1000100000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=380
      ("1001000000100010", '0', '1', "01", "010", "010", "000", '0', '-', "00"), -- i=381
      ("1001100000100010", '1', '1', "01", "010", "010", "000", '0', '-', "00"), -- i=382
      ("1001100000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=383
      ("1010000000100010", '0', '1', "10", "010", "010", "000", '0', '-', "00"), -- i=384
      ("1010100000100010", '1', '1', "10", "010", "010", "000", '0', '-', "00"), -- i=385
      ("1010100000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=386
      ("1011000000100010", '0', '1', "11", "010", "010", "000", '0', '-', "00"), -- i=387
      ("1011100000100010", '1', '1', "11", "010", "010", "000", '0', '-', "00"), -- i=388
      ("1011100000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=389
      ("0101000000100000", '0', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=390
      ("0101100000100000", '1', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=391
      ("0101100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=392
      ("0100000000100000", '0', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=393
      ("0100100000100000", '1', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=394
      ("0100100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=395
      ("0000000000101000", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=396
      ("0000100000101000", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=397
      ("0000100000101000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=398
      ("1000000000100011", '0', '1', "00", "010", "011", "000", '0', '-', "00"), -- i=399
      ("1000100000100011", '1', '1', "00", "010", "011", "000", '0', '-', "00"), -- i=400
      ("1000100000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=401
      ("1001000000100011", '0', '1', "01", "010", "011", "000", '0', '-', "00"), -- i=402
      ("1001100000100011", '1', '1', "01", "010", "011", "000", '0', '-', "00"), -- i=403
      ("1001100000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=404
      ("1010000000100011", '0', '1', "10", "010", "011", "000", '0', '-', "00"), -- i=405
      ("1010100000100011", '1', '1', "10", "010", "011", "000", '0', '-', "00"), -- i=406
      ("1010100000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=407
      ("1011000000100011", '0', '1', "11", "010", "011", "000", '0', '-', "00"), -- i=408
      ("1011100000100011", '1', '1', "11", "010", "011", "000", '0', '-', "00"), -- i=409
      ("1011100000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=410
      ("0101000000100000", '0', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=411
      ("0101100000100000", '1', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=412
      ("0101100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=413
      ("0100000000100000", '0', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=414
      ("0100100000100000", '1', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=415
      ("0100100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=416
      ("0000000001001001", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=417
      ("0000100001001001", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=418
      ("0000100001001001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=419
      ("1000000000100100", '0', '1', "00", "010", "100", "000", '0', '-', "00"), -- i=420
      ("1000100000100100", '1', '1', "00", "010", "100", "000", '0', '-', "00"), -- i=421
      ("1000100000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=422
      ("1001000000100100", '0', '1', "01", "010", "100", "000", '0', '-', "00"), -- i=423
      ("1001100000100100", '1', '1', "01", "010", "100", "000", '0', '-', "00"), -- i=424
      ("1001100000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=425
      ("1010000000100100", '0', '1', "10", "010", "100", "000", '0', '-', "00"), -- i=426
      ("1010100000100100", '1', '1', "10", "010", "100", "000", '0', '-', "00"), -- i=427
      ("1010100000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=428
      ("1011000000100100", '0', '1', "11", "010", "100", "000", '0', '-', "00"), -- i=429
      ("1011100000100100", '1', '1', "11", "010", "100", "000", '0', '-', "00"), -- i=430
      ("1011100000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=431
      ("0101000000100000", '0', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=432
      ("0101100000100000", '1', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=433
      ("0101100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=434
      ("0100000000100000", '0', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=435
      ("0100100000100000", '1', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=436
      ("0100100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=437
      ("0000000001000011", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=438
      ("0000100001000011", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=439
      ("0000100001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=440
      ("1000000000100101", '0', '1', "00", "010", "101", "000", '0', '-', "00"), -- i=441
      ("1000100000100101", '1', '1', "00", "010", "101", "000", '0', '-', "00"), -- i=442
      ("1000100000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=443
      ("1001000000100101", '0', '1', "01", "010", "101", "000", '0', '-', "00"), -- i=444
      ("1001100000100101", '1', '1', "01", "010", "101", "000", '0', '-', "00"), -- i=445
      ("1001100000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=446
      ("1010000000100101", '0', '1', "10", "010", "101", "000", '0', '-', "00"), -- i=447
      ("1010100000100101", '1', '1', "10", "010", "101", "000", '0', '-', "00"), -- i=448
      ("1010100000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=449
      ("1011000000100101", '0', '1', "11", "010", "101", "000", '0', '-', "00"), -- i=450
      ("1011100000100101", '1', '1', "11", "010", "101", "000", '0', '-', "00"), -- i=451
      ("1011100000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=452
      ("0101000000100000", '0', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=453
      ("0101100000100000", '1', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=454
      ("0101100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=455
      ("0100000000100000", '0', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=456
      ("0100100000100000", '1', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=457
      ("0100100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=458
      ("0000000010010011", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=459
      ("0000100010010011", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=460
      ("0000100010010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=461
      ("1000000000100110", '0', '1', "00", "010", "110", "000", '0', '-', "00"), -- i=462
      ("1000100000100110", '1', '1', "00", "010", "110", "000", '0', '-', "00"), -- i=463
      ("1000100000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=464
      ("1001000000100110", '0', '1', "01", "010", "110", "000", '0', '-', "00"), -- i=465
      ("1001100000100110", '1', '1', "01", "010", "110", "000", '0', '-', "00"), -- i=466
      ("1001100000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=467
      ("1010000000100110", '0', '1', "10", "010", "110", "000", '0', '-', "00"), -- i=468
      ("1010100000100110", '1', '1', "10", "010", "110", "000", '0', '-', "00"), -- i=469
      ("1010100000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=470
      ("1011000000100110", '0', '1', "11", "010", "110", "000", '0', '-', "00"), -- i=471
      ("1011100000100110", '1', '1', "11", "010", "110", "000", '0', '-', "00"), -- i=472
      ("1011100000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=473
      ("0101000000100000", '0', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=474
      ("0101100000100000", '1', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=475
      ("0101100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=476
      ("0100000000100000", '0', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=477
      ("0100100000100000", '1', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=478
      ("0100100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=479
      ("0000000010010111", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=480
      ("0000100010010111", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=481
      ("0000100010010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=482
      ("1000000000100111", '0', '1', "00", "010", "111", "000", '0', '-', "00"), -- i=483
      ("1000100000100111", '1', '1', "00", "010", "111", "000", '0', '-', "00"), -- i=484
      ("1000100000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=485
      ("1001000000100111", '0', '1', "01", "010", "111", "000", '0', '-', "00"), -- i=486
      ("1001100000100111", '1', '1', "01", "010", "111", "000", '0', '-', "00"), -- i=487
      ("1001100000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=488
      ("1010000000100111", '0', '1', "10", "010", "111", "000", '0', '-', "00"), -- i=489
      ("1010100000100111", '1', '1', "10", "010", "111", "000", '0', '-', "00"), -- i=490
      ("1010100000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=491
      ("1011000000100111", '0', '1', "11", "010", "111", "000", '0', '-', "00"), -- i=492
      ("1011100000100111", '1', '1', "11", "010", "111", "000", '0', '-', "00"), -- i=493
      ("1011100000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=494
      ("0101000000100000", '0', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=495
      ("0101100000100000", '1', '1', "--", "010", "---", "000", '0', '1', "01"), -- i=496
      ("0101100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=497
      ("0100000000100000", '0', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=498
      ("0100100000100000", '1', '0', "--", "010", "000", "---", '1', '-', "--"), -- i=499
      ("0100100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=500
      ("0000000000100100", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=501
      ("0000100000100100", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=502
      ("0000100000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=503
      ("1000000000110000", '0', '1', "00", "011", "000", "000", '0', '-', "00"), -- i=504
      ("1000100000110000", '1', '1', "00", "011", "000", "000", '0', '-', "00"), -- i=505
      ("1000100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=506
      ("1001000000110000", '0', '1', "01", "011", "000", "000", '0', '-', "00"), -- i=507
      ("1001100000110000", '1', '1', "01", "011", "000", "000", '0', '-', "00"), -- i=508
      ("1001100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=509
      ("1010000000110000", '0', '1', "10", "011", "000", "000", '0', '-', "00"), -- i=510
      ("1010100000110000", '1', '1', "10", "011", "000", "000", '0', '-', "00"), -- i=511
      ("1010100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=512
      ("1011000000110000", '0', '1', "11", "011", "000", "000", '0', '-', "00"), -- i=513
      ("1011100000110000", '1', '1', "11", "011", "000", "000", '0', '-', "00"), -- i=514
      ("1011100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=515
      ("0101000000110000", '0', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=516
      ("0101100000110000", '1', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=517
      ("0101100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=518
      ("0100000000110000", '0', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=519
      ("0100100000110000", '1', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=520
      ("0100100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=521
      ("0000000001001000", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=522
      ("0000100001001000", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=523
      ("0000100001001000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=524
      ("1000000000110001", '0', '1', "00", "011", "001", "000", '0', '-', "00"), -- i=525
      ("1000100000110001", '1', '1', "00", "011", "001", "000", '0', '-', "00"), -- i=526
      ("1000100000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=527
      ("1001000000110001", '0', '1', "01", "011", "001", "000", '0', '-', "00"), -- i=528
      ("1001100000110001", '1', '1', "01", "011", "001", "000", '0', '-', "00"), -- i=529
      ("1001100000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=530
      ("1010000000110001", '0', '1', "10", "011", "001", "000", '0', '-', "00"), -- i=531
      ("1010100000110001", '1', '1', "10", "011", "001", "000", '0', '-', "00"), -- i=532
      ("1010100000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=533
      ("1011000000110001", '0', '1', "11", "011", "001", "000", '0', '-', "00"), -- i=534
      ("1011100000110001", '1', '1', "11", "011", "001", "000", '0', '-', "00"), -- i=535
      ("1011100000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=536
      ("0101000000110000", '0', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=537
      ("0101100000110000", '1', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=538
      ("0101100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=539
      ("0100000000110000", '0', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=540
      ("0100100000110000", '1', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=541
      ("0100100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=542
      ("0000000010100110", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=543
      ("0000100010100110", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=544
      ("0000100010100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=545
      ("1000000000110010", '0', '1', "00", "011", "010", "000", '0', '-', "00"), -- i=546
      ("1000100000110010", '1', '1', "00", "011", "010", "000", '0', '-', "00"), -- i=547
      ("1000100000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=548
      ("1001000000110010", '0', '1', "01", "011", "010", "000", '0', '-', "00"), -- i=549
      ("1001100000110010", '1', '1', "01", "011", "010", "000", '0', '-', "00"), -- i=550
      ("1001100000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=551
      ("1010000000110010", '0', '1', "10", "011", "010", "000", '0', '-', "00"), -- i=552
      ("1010100000110010", '1', '1', "10", "011", "010", "000", '0', '-', "00"), -- i=553
      ("1010100000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=554
      ("1011000000110010", '0', '1', "11", "011", "010", "000", '0', '-', "00"), -- i=555
      ("1011100000110010", '1', '1', "11", "011", "010", "000", '0', '-', "00"), -- i=556
      ("1011100000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=557
      ("0101000000110000", '0', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=558
      ("0101100000110000", '1', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=559
      ("0101100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=560
      ("0100000000110000", '0', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=561
      ("0100100000110000", '1', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=562
      ("0100100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=563
      ("0000000010111101", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=564
      ("0000100010111101", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=565
      ("0000100010111101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=566
      ("1000000000110011", '0', '1', "00", "011", "011", "000", '0', '-', "00"), -- i=567
      ("1000100000110011", '1', '1', "00", "011", "011", "000", '0', '-', "00"), -- i=568
      ("1000100000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=569
      ("1001000000110011", '0', '1', "01", "011", "011", "000", '0', '-', "00"), -- i=570
      ("1001100000110011", '1', '1', "01", "011", "011", "000", '0', '-', "00"), -- i=571
      ("1001100000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=572
      ("1010000000110011", '0', '1', "10", "011", "011", "000", '0', '-', "00"), -- i=573
      ("1010100000110011", '1', '1', "10", "011", "011", "000", '0', '-', "00"), -- i=574
      ("1010100000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=575
      ("1011000000110011", '0', '1', "11", "011", "011", "000", '0', '-', "00"), -- i=576
      ("1011100000110011", '1', '1', "11", "011", "011", "000", '0', '-', "00"), -- i=577
      ("1011100000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=578
      ("0101000000110000", '0', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=579
      ("0101100000110000", '1', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=580
      ("0101100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=581
      ("0100000000110000", '0', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=582
      ("0100100000110000", '1', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=583
      ("0100100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=584
      ("0000000001011110", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=585
      ("0000100001011110", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=586
      ("0000100001011110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=587
      ("1000000000110100", '0', '1', "00", "011", "100", "000", '0', '-', "00"), -- i=588
      ("1000100000110100", '1', '1', "00", "011", "100", "000", '0', '-', "00"), -- i=589
      ("1000100000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=590
      ("1001000000110100", '0', '1', "01", "011", "100", "000", '0', '-', "00"), -- i=591
      ("1001100000110100", '1', '1', "01", "011", "100", "000", '0', '-', "00"), -- i=592
      ("1001100000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=593
      ("1010000000110100", '0', '1', "10", "011", "100", "000", '0', '-', "00"), -- i=594
      ("1010100000110100", '1', '1', "10", "011", "100", "000", '0', '-', "00"), -- i=595
      ("1010100000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=596
      ("1011000000110100", '0', '1', "11", "011", "100", "000", '0', '-', "00"), -- i=597
      ("1011100000110100", '1', '1', "11", "011", "100", "000", '0', '-', "00"), -- i=598
      ("1011100000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=599
      ("0101000000110000", '0', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=600
      ("0101100000110000", '1', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=601
      ("0101100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=602
      ("0100000000110000", '0', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=603
      ("0100100000110000", '1', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=604
      ("0100100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=605
      ("0000000011110110", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=606
      ("0000100011110110", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=607
      ("0000100011110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=608
      ("1000000000110101", '0', '1', "00", "011", "101", "000", '0', '-', "00"), -- i=609
      ("1000100000110101", '1', '1', "00", "011", "101", "000", '0', '-', "00"), -- i=610
      ("1000100000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=611
      ("1001000000110101", '0', '1', "01", "011", "101", "000", '0', '-', "00"), -- i=612
      ("1001100000110101", '1', '1', "01", "011", "101", "000", '0', '-', "00"), -- i=613
      ("1001100000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=614
      ("1010000000110101", '0', '1', "10", "011", "101", "000", '0', '-', "00"), -- i=615
      ("1010100000110101", '1', '1', "10", "011", "101", "000", '0', '-', "00"), -- i=616
      ("1010100000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=617
      ("1011000000110101", '0', '1', "11", "011", "101", "000", '0', '-', "00"), -- i=618
      ("1011100000110101", '1', '1', "11", "011", "101", "000", '0', '-', "00"), -- i=619
      ("1011100000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=620
      ("0101000000110000", '0', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=621
      ("0101100000110000", '1', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=622
      ("0101100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=623
      ("0100000000110000", '0', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=624
      ("0100100000110000", '1', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=625
      ("0100100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=626
      ("0000000001000000", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=627
      ("0000100001000000", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=628
      ("0000100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=629
      ("1000000000110110", '0', '1', "00", "011", "110", "000", '0', '-', "00"), -- i=630
      ("1000100000110110", '1', '1', "00", "011", "110", "000", '0', '-', "00"), -- i=631
      ("1000100000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=632
      ("1001000000110110", '0', '1', "01", "011", "110", "000", '0', '-', "00"), -- i=633
      ("1001100000110110", '1', '1', "01", "011", "110", "000", '0', '-', "00"), -- i=634
      ("1001100000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=635
      ("1010000000110110", '0', '1', "10", "011", "110", "000", '0', '-', "00"), -- i=636
      ("1010100000110110", '1', '1', "10", "011", "110", "000", '0', '-', "00"), -- i=637
      ("1010100000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=638
      ("1011000000110110", '0', '1', "11", "011", "110", "000", '0', '-', "00"), -- i=639
      ("1011100000110110", '1', '1', "11", "011", "110", "000", '0', '-', "00"), -- i=640
      ("1011100000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=641
      ("0101000000110000", '0', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=642
      ("0101100000110000", '1', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=643
      ("0101100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=644
      ("0100000000110000", '0', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=645
      ("0100100000110000", '1', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=646
      ("0100100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=647
      ("0000000000111001", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=648
      ("0000100000111001", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=649
      ("0000100000111001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=650
      ("1000000000110111", '0', '1', "00", "011", "111", "000", '0', '-', "00"), -- i=651
      ("1000100000110111", '1', '1', "00", "011", "111", "000", '0', '-', "00"), -- i=652
      ("1000100000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=653
      ("1001000000110111", '0', '1', "01", "011", "111", "000", '0', '-', "00"), -- i=654
      ("1001100000110111", '1', '1', "01", "011", "111", "000", '0', '-', "00"), -- i=655
      ("1001100000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=656
      ("1010000000110111", '0', '1', "10", "011", "111", "000", '0', '-', "00"), -- i=657
      ("1010100000110111", '1', '1', "10", "011", "111", "000", '0', '-', "00"), -- i=658
      ("1010100000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=659
      ("1011000000110111", '0', '1', "11", "011", "111", "000", '0', '-', "00"), -- i=660
      ("1011100000110111", '1', '1', "11", "011", "111", "000", '0', '-', "00"), -- i=661
      ("1011100000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=662
      ("0101000000110000", '0', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=663
      ("0101100000110000", '1', '1', "--", "011", "---", "000", '0', '1', "01"), -- i=664
      ("0101100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=665
      ("0100000000110000", '0', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=666
      ("0100100000110000", '1', '0', "--", "011", "000", "---", '1', '-', "--"), -- i=667
      ("0100100000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=668
      ("0000000010101000", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=669
      ("0000100010101000", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=670
      ("0000100010101000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=671
      ("1000000001000000", '0', '1', "00", "100", "000", "000", '0', '-', "00"), -- i=672
      ("1000100001000000", '1', '1', "00", "100", "000", "000", '0', '-', "00"), -- i=673
      ("1000100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=674
      ("1001000001000000", '0', '1', "01", "100", "000", "000", '0', '-', "00"), -- i=675
      ("1001100001000000", '1', '1', "01", "100", "000", "000", '0', '-', "00"), -- i=676
      ("1001100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=677
      ("1010000001000000", '0', '1', "10", "100", "000", "000", '0', '-', "00"), -- i=678
      ("1010100001000000", '1', '1', "10", "100", "000", "000", '0', '-', "00"), -- i=679
      ("1010100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=680
      ("1011000001000000", '0', '1', "11", "100", "000", "000", '0', '-', "00"), -- i=681
      ("1011100001000000", '1', '1', "11", "100", "000", "000", '0', '-', "00"), -- i=682
      ("1011100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=683
      ("0101000001000000", '0', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=684
      ("0101100001000000", '1', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=685
      ("0101100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=686
      ("0100000001000000", '0', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=687
      ("0100100001000000", '1', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=688
      ("0100100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=689
      ("0000000001100000", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=690
      ("0000100001100000", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=691
      ("0000100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=692
      ("1000000001000001", '0', '1', "00", "100", "001", "000", '0', '-', "00"), -- i=693
      ("1000100001000001", '1', '1', "00", "100", "001", "000", '0', '-', "00"), -- i=694
      ("1000100001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=695
      ("1001000001000001", '0', '1', "01", "100", "001", "000", '0', '-', "00"), -- i=696
      ("1001100001000001", '1', '1', "01", "100", "001", "000", '0', '-', "00"), -- i=697
      ("1001100001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=698
      ("1010000001000001", '0', '1', "10", "100", "001", "000", '0', '-', "00"), -- i=699
      ("1010100001000001", '1', '1', "10", "100", "001", "000", '0', '-', "00"), -- i=700
      ("1010100001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=701
      ("1011000001000001", '0', '1', "11", "100", "001", "000", '0', '-', "00"), -- i=702
      ("1011100001000001", '1', '1', "11", "100", "001", "000", '0', '-', "00"), -- i=703
      ("1011100001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=704
      ("0101000001000000", '0', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=705
      ("0101100001000000", '1', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=706
      ("0101100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=707
      ("0100000001000000", '0', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=708
      ("0100100001000000", '1', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=709
      ("0100100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=710
      ("0000000000010101", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=711
      ("0000100000010101", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=712
      ("0000100000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=713
      ("1000000001000010", '0', '1', "00", "100", "010", "000", '0', '-', "00"), -- i=714
      ("1000100001000010", '1', '1', "00", "100", "010", "000", '0', '-', "00"), -- i=715
      ("1000100001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=716
      ("1001000001000010", '0', '1', "01", "100", "010", "000", '0', '-', "00"), -- i=717
      ("1001100001000010", '1', '1', "01", "100", "010", "000", '0', '-', "00"), -- i=718
      ("1001100001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=719
      ("1010000001000010", '0', '1', "10", "100", "010", "000", '0', '-', "00"), -- i=720
      ("1010100001000010", '1', '1', "10", "100", "010", "000", '0', '-', "00"), -- i=721
      ("1010100001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=722
      ("1011000001000010", '0', '1', "11", "100", "010", "000", '0', '-', "00"), -- i=723
      ("1011100001000010", '1', '1', "11", "100", "010", "000", '0', '-', "00"), -- i=724
      ("1011100001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=725
      ("0101000001000000", '0', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=726
      ("0101100001000000", '1', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=727
      ("0101100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=728
      ("0100000001000000", '0', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=729
      ("0100100001000000", '1', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=730
      ("0100100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=731
      ("0000000000111000", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=732
      ("0000100000111000", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=733
      ("0000100000111000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=734
      ("1000000001000011", '0', '1', "00", "100", "011", "000", '0', '-', "00"), -- i=735
      ("1000100001000011", '1', '1', "00", "100", "011", "000", '0', '-', "00"), -- i=736
      ("1000100001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=737
      ("1001000001000011", '0', '1', "01", "100", "011", "000", '0', '-', "00"), -- i=738
      ("1001100001000011", '1', '1', "01", "100", "011", "000", '0', '-', "00"), -- i=739
      ("1001100001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=740
      ("1010000001000011", '0', '1', "10", "100", "011", "000", '0', '-', "00"), -- i=741
      ("1010100001000011", '1', '1', "10", "100", "011", "000", '0', '-', "00"), -- i=742
      ("1010100001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=743
      ("1011000001000011", '0', '1', "11", "100", "011", "000", '0', '-', "00"), -- i=744
      ("1011100001000011", '1', '1', "11", "100", "011", "000", '0', '-', "00"), -- i=745
      ("1011100001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=746
      ("0101000001000000", '0', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=747
      ("0101100001000000", '1', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=748
      ("0101100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=749
      ("0100000001000000", '0', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=750
      ("0100100001000000", '1', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=751
      ("0100100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=752
      ("0000000000100000", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=753
      ("0000100000100000", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=754
      ("0000100000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=755
      ("1000000001000100", '0', '1', "00", "100", "100", "000", '0', '-', "00"), -- i=756
      ("1000100001000100", '1', '1', "00", "100", "100", "000", '0', '-', "00"), -- i=757
      ("1000100001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=758
      ("1001000001000100", '0', '1', "01", "100", "100", "000", '0', '-', "00"), -- i=759
      ("1001100001000100", '1', '1', "01", "100", "100", "000", '0', '-', "00"), -- i=760
      ("1001100001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=761
      ("1010000001000100", '0', '1', "10", "100", "100", "000", '0', '-', "00"), -- i=762
      ("1010100001000100", '1', '1', "10", "100", "100", "000", '0', '-', "00"), -- i=763
      ("1010100001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=764
      ("1011000001000100", '0', '1', "11", "100", "100", "000", '0', '-', "00"), -- i=765
      ("1011100001000100", '1', '1', "11", "100", "100", "000", '0', '-', "00"), -- i=766
      ("1011100001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=767
      ("0101000001000000", '0', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=768
      ("0101100001000000", '1', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=769
      ("0101100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=770
      ("0100000001000000", '0', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=771
      ("0100100001000000", '1', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=772
      ("0100100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=773
      ("0000000010111010", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=774
      ("0000100010111010", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=775
      ("0000100010111010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=776
      ("1000000001000101", '0', '1', "00", "100", "101", "000", '0', '-', "00"), -- i=777
      ("1000100001000101", '1', '1', "00", "100", "101", "000", '0', '-', "00"), -- i=778
      ("1000100001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=779
      ("1001000001000101", '0', '1', "01", "100", "101", "000", '0', '-', "00"), -- i=780
      ("1001100001000101", '1', '1', "01", "100", "101", "000", '0', '-', "00"), -- i=781
      ("1001100001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=782
      ("1010000001000101", '0', '1', "10", "100", "101", "000", '0', '-', "00"), -- i=783
      ("1010100001000101", '1', '1', "10", "100", "101", "000", '0', '-', "00"), -- i=784
      ("1010100001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=785
      ("1011000001000101", '0', '1', "11", "100", "101", "000", '0', '-', "00"), -- i=786
      ("1011100001000101", '1', '1', "11", "100", "101", "000", '0', '-', "00"), -- i=787
      ("1011100001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=788
      ("0101000001000000", '0', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=789
      ("0101100001000000", '1', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=790
      ("0101100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=791
      ("0100000001000000", '0', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=792
      ("0100100001000000", '1', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=793
      ("0100100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=794
      ("0000000001110001", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=795
      ("0000100001110001", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=796
      ("0000100001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=797
      ("1000000001000110", '0', '1', "00", "100", "110", "000", '0', '-', "00"), -- i=798
      ("1000100001000110", '1', '1', "00", "100", "110", "000", '0', '-', "00"), -- i=799
      ("1000100001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=800
      ("1001000001000110", '0', '1', "01", "100", "110", "000", '0', '-', "00"), -- i=801
      ("1001100001000110", '1', '1', "01", "100", "110", "000", '0', '-', "00"), -- i=802
      ("1001100001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=803
      ("1010000001000110", '0', '1', "10", "100", "110", "000", '0', '-', "00"), -- i=804
      ("1010100001000110", '1', '1', "10", "100", "110", "000", '0', '-', "00"), -- i=805
      ("1010100001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=806
      ("1011000001000110", '0', '1', "11", "100", "110", "000", '0', '-', "00"), -- i=807
      ("1011100001000110", '1', '1', "11", "100", "110", "000", '0', '-', "00"), -- i=808
      ("1011100001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=809
      ("0101000001000000", '0', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=810
      ("0101100001000000", '1', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=811
      ("0101100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=812
      ("0100000001000000", '0', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=813
      ("0100100001000000", '1', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=814
      ("0100100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=815
      ("0000000010011010", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=816
      ("0000100010011010", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=817
      ("0000100010011010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=818
      ("1000000001000111", '0', '1', "00", "100", "111", "000", '0', '-', "00"), -- i=819
      ("1000100001000111", '1', '1', "00", "100", "111", "000", '0', '-', "00"), -- i=820
      ("1000100001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=821
      ("1001000001000111", '0', '1', "01", "100", "111", "000", '0', '-', "00"), -- i=822
      ("1001100001000111", '1', '1', "01", "100", "111", "000", '0', '-', "00"), -- i=823
      ("1001100001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=824
      ("1010000001000111", '0', '1', "10", "100", "111", "000", '0', '-', "00"), -- i=825
      ("1010100001000111", '1', '1', "10", "100", "111", "000", '0', '-', "00"), -- i=826
      ("1010100001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=827
      ("1011000001000111", '0', '1', "11", "100", "111", "000", '0', '-', "00"), -- i=828
      ("1011100001000111", '1', '1', "11", "100", "111", "000", '0', '-', "00"), -- i=829
      ("1011100001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=830
      ("0101000001000000", '0', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=831
      ("0101100001000000", '1', '1', "--", "100", "---", "000", '0', '1', "01"), -- i=832
      ("0101100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=833
      ("0100000001000000", '0', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=834
      ("0100100001000000", '1', '0', "--", "100", "000", "---", '1', '-', "--"), -- i=835
      ("0100100001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=836
      ("0000000001010010", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=837
      ("0000100001010010", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=838
      ("0000100001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=839
      ("1000000001010000", '0', '1', "00", "101", "000", "000", '0', '-', "00"), -- i=840
      ("1000100001010000", '1', '1', "00", "101", "000", "000", '0', '-', "00"), -- i=841
      ("1000100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=842
      ("1001000001010000", '0', '1', "01", "101", "000", "000", '0', '-', "00"), -- i=843
      ("1001100001010000", '1', '1', "01", "101", "000", "000", '0', '-', "00"), -- i=844
      ("1001100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=845
      ("1010000001010000", '0', '1', "10", "101", "000", "000", '0', '-', "00"), -- i=846
      ("1010100001010000", '1', '1', "10", "101", "000", "000", '0', '-', "00"), -- i=847
      ("1010100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=848
      ("1011000001010000", '0', '1', "11", "101", "000", "000", '0', '-', "00"), -- i=849
      ("1011100001010000", '1', '1', "11", "101", "000", "000", '0', '-', "00"), -- i=850
      ("1011100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=851
      ("0101000001010000", '0', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=852
      ("0101100001010000", '1', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=853
      ("0101100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=854
      ("0100000001010000", '0', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=855
      ("0100100001010000", '1', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=856
      ("0100100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=857
      ("0000000001111100", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=858
      ("0000100001111100", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=859
      ("0000100001111100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=860
      ("1000000001010001", '0', '1', "00", "101", "001", "000", '0', '-', "00"), -- i=861
      ("1000100001010001", '1', '1', "00", "101", "001", "000", '0', '-', "00"), -- i=862
      ("1000100001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=863
      ("1001000001010001", '0', '1', "01", "101", "001", "000", '0', '-', "00"), -- i=864
      ("1001100001010001", '1', '1', "01", "101", "001", "000", '0', '-', "00"), -- i=865
      ("1001100001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=866
      ("1010000001010001", '0', '1', "10", "101", "001", "000", '0', '-', "00"), -- i=867
      ("1010100001010001", '1', '1', "10", "101", "001", "000", '0', '-', "00"), -- i=868
      ("1010100001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=869
      ("1011000001010001", '0', '1', "11", "101", "001", "000", '0', '-', "00"), -- i=870
      ("1011100001010001", '1', '1', "11", "101", "001", "000", '0', '-', "00"), -- i=871
      ("1011100001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=872
      ("0101000001010000", '0', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=873
      ("0101100001010000", '1', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=874
      ("0101100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=875
      ("0100000001010000", '0', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=876
      ("0100100001010000", '1', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=877
      ("0100100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=878
      ("0000000000101110", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=879
      ("0000100000101110", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=880
      ("0000100000101110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=881
      ("1000000001010010", '0', '1', "00", "101", "010", "000", '0', '-', "00"), -- i=882
      ("1000100001010010", '1', '1', "00", "101", "010", "000", '0', '-', "00"), -- i=883
      ("1000100001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=884
      ("1001000001010010", '0', '1', "01", "101", "010", "000", '0', '-', "00"), -- i=885
      ("1001100001010010", '1', '1', "01", "101", "010", "000", '0', '-', "00"), -- i=886
      ("1001100001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=887
      ("1010000001010010", '0', '1', "10", "101", "010", "000", '0', '-', "00"), -- i=888
      ("1010100001010010", '1', '1', "10", "101", "010", "000", '0', '-', "00"), -- i=889
      ("1010100001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=890
      ("1011000001010010", '0', '1', "11", "101", "010", "000", '0', '-', "00"), -- i=891
      ("1011100001010010", '1', '1', "11", "101", "010", "000", '0', '-', "00"), -- i=892
      ("1011100001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=893
      ("0101000001010000", '0', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=894
      ("0101100001010000", '1', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=895
      ("0101100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=896
      ("0100000001010000", '0', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=897
      ("0100100001010000", '1', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=898
      ("0100100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=899
      ("0000000011000011", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=900
      ("0000100011000011", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=901
      ("0000100011000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=902
      ("1000000001010011", '0', '1', "00", "101", "011", "000", '0', '-', "00"), -- i=903
      ("1000100001010011", '1', '1', "00", "101", "011", "000", '0', '-', "00"), -- i=904
      ("1000100001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=905
      ("1001000001010011", '0', '1', "01", "101", "011", "000", '0', '-', "00"), -- i=906
      ("1001100001010011", '1', '1', "01", "101", "011", "000", '0', '-', "00"), -- i=907
      ("1001100001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=908
      ("1010000001010011", '0', '1', "10", "101", "011", "000", '0', '-', "00"), -- i=909
      ("1010100001010011", '1', '1', "10", "101", "011", "000", '0', '-', "00"), -- i=910
      ("1010100001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=911
      ("1011000001010011", '0', '1', "11", "101", "011", "000", '0', '-', "00"), -- i=912
      ("1011100001010011", '1', '1', "11", "101", "011", "000", '0', '-', "00"), -- i=913
      ("1011100001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=914
      ("0101000001010000", '0', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=915
      ("0101100001010000", '1', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=916
      ("0101100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=917
      ("0100000001010000", '0', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=918
      ("0100100001010000", '1', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=919
      ("0100100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=920
      ("0000000010010001", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=921
      ("0000100010010001", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=922
      ("0000100010010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=923
      ("1000000001010100", '0', '1', "00", "101", "100", "000", '0', '-', "00"), -- i=924
      ("1000100001010100", '1', '1', "00", "101", "100", "000", '0', '-', "00"), -- i=925
      ("1000100001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=926
      ("1001000001010100", '0', '1', "01", "101", "100", "000", '0', '-', "00"), -- i=927
      ("1001100001010100", '1', '1', "01", "101", "100", "000", '0', '-', "00"), -- i=928
      ("1001100001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=929
      ("1010000001010100", '0', '1', "10", "101", "100", "000", '0', '-', "00"), -- i=930
      ("1010100001010100", '1', '1', "10", "101", "100", "000", '0', '-', "00"), -- i=931
      ("1010100001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=932
      ("1011000001010100", '0', '1', "11", "101", "100", "000", '0', '-', "00"), -- i=933
      ("1011100001010100", '1', '1', "11", "101", "100", "000", '0', '-', "00"), -- i=934
      ("1011100001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=935
      ("0101000001010000", '0', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=936
      ("0101100001010000", '1', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=937
      ("0101100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=938
      ("0100000001010000", '0', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=939
      ("0100100001010000", '1', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=940
      ("0100100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=941
      ("0000000011010010", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=942
      ("0000100011010010", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=943
      ("0000100011010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=944
      ("1000000001010101", '0', '1', "00", "101", "101", "000", '0', '-', "00"), -- i=945
      ("1000100001010101", '1', '1', "00", "101", "101", "000", '0', '-', "00"), -- i=946
      ("1000100001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=947
      ("1001000001010101", '0', '1', "01", "101", "101", "000", '0', '-', "00"), -- i=948
      ("1001100001010101", '1', '1', "01", "101", "101", "000", '0', '-', "00"), -- i=949
      ("1001100001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=950
      ("1010000001010101", '0', '1', "10", "101", "101", "000", '0', '-', "00"), -- i=951
      ("1010100001010101", '1', '1', "10", "101", "101", "000", '0', '-', "00"), -- i=952
      ("1010100001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=953
      ("1011000001010101", '0', '1', "11", "101", "101", "000", '0', '-', "00"), -- i=954
      ("1011100001010101", '1', '1', "11", "101", "101", "000", '0', '-', "00"), -- i=955
      ("1011100001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=956
      ("0101000001010000", '0', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=957
      ("0101100001010000", '1', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=958
      ("0101100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=959
      ("0100000001010000", '0', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=960
      ("0100100001010000", '1', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=961
      ("0100100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=962
      ("0000000010110011", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=963
      ("0000100010110011", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=964
      ("0000100010110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=965
      ("1000000001010110", '0', '1', "00", "101", "110", "000", '0', '-', "00"), -- i=966
      ("1000100001010110", '1', '1', "00", "101", "110", "000", '0', '-', "00"), -- i=967
      ("1000100001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=968
      ("1001000001010110", '0', '1', "01", "101", "110", "000", '0', '-', "00"), -- i=969
      ("1001100001010110", '1', '1', "01", "101", "110", "000", '0', '-', "00"), -- i=970
      ("1001100001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=971
      ("1010000001010110", '0', '1', "10", "101", "110", "000", '0', '-', "00"), -- i=972
      ("1010100001010110", '1', '1', "10", "101", "110", "000", '0', '-', "00"), -- i=973
      ("1010100001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=974
      ("1011000001010110", '0', '1', "11", "101", "110", "000", '0', '-', "00"), -- i=975
      ("1011100001010110", '1', '1', "11", "101", "110", "000", '0', '-', "00"), -- i=976
      ("1011100001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=977
      ("0101000001010000", '0', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=978
      ("0101100001010000", '1', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=979
      ("0101100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=980
      ("0100000001010000", '0', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=981
      ("0100100001010000", '1', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=982
      ("0100100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=983
      ("0000000001010110", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=984
      ("0000100001010110", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=985
      ("0000100001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=986
      ("1000000001010111", '0', '1', "00", "101", "111", "000", '0', '-', "00"), -- i=987
      ("1000100001010111", '1', '1', "00", "101", "111", "000", '0', '-', "00"), -- i=988
      ("1000100001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=989
      ("1001000001010111", '0', '1', "01", "101", "111", "000", '0', '-', "00"), -- i=990
      ("1001100001010111", '1', '1', "01", "101", "111", "000", '0', '-', "00"), -- i=991
      ("1001100001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=992
      ("1010000001010111", '0', '1', "10", "101", "111", "000", '0', '-', "00"), -- i=993
      ("1010100001010111", '1', '1', "10", "101", "111", "000", '0', '-', "00"), -- i=994
      ("1010100001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=995
      ("1011000001010111", '0', '1', "11", "101", "111", "000", '0', '-', "00"), -- i=996
      ("1011100001010111", '1', '1', "11", "101", "111", "000", '0', '-', "00"), -- i=997
      ("1011100001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=998
      ("0101000001010000", '0', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=999
      ("0101100001010000", '1', '1', "--", "101", "---", "000", '0', '1', "01"), -- i=1000
      ("0101100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1001
      ("0100000001010000", '0', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=1002
      ("0100100001010000", '1', '0', "--", "101", "000", "---", '1', '-', "--"), -- i=1003
      ("0100100001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1004
      ("0000000010101110", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1005
      ("0000100010101110", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1006
      ("0000100010101110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1007
      ("1000000001100000", '0', '1', "00", "110", "000", "000", '0', '-', "00"), -- i=1008
      ("1000100001100000", '1', '1', "00", "110", "000", "000", '0', '-', "00"), -- i=1009
      ("1000100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1010
      ("1001000001100000", '0', '1', "01", "110", "000", "000", '0', '-', "00"), -- i=1011
      ("1001100001100000", '1', '1', "01", "110", "000", "000", '0', '-', "00"), -- i=1012
      ("1001100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1013
      ("1010000001100000", '0', '1', "10", "110", "000", "000", '0', '-', "00"), -- i=1014
      ("1010100001100000", '1', '1', "10", "110", "000", "000", '0', '-', "00"), -- i=1015
      ("1010100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1016
      ("1011000001100000", '0', '1', "11", "110", "000", "000", '0', '-', "00"), -- i=1017
      ("1011100001100000", '1', '1', "11", "110", "000", "000", '0', '-', "00"), -- i=1018
      ("1011100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1019
      ("0101000001100000", '0', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1020
      ("0101100001100000", '1', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1021
      ("0101100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1022
      ("0100000001100000", '0', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1023
      ("0100100001100000", '1', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1024
      ("0100100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1025
      ("0000000010111011", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1026
      ("0000100010111011", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1027
      ("0000100010111011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1028
      ("1000000001100001", '0', '1', "00", "110", "001", "000", '0', '-', "00"), -- i=1029
      ("1000100001100001", '1', '1', "00", "110", "001", "000", '0', '-', "00"), -- i=1030
      ("1000100001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1031
      ("1001000001100001", '0', '1', "01", "110", "001", "000", '0', '-', "00"), -- i=1032
      ("1001100001100001", '1', '1', "01", "110", "001", "000", '0', '-', "00"), -- i=1033
      ("1001100001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1034
      ("1010000001100001", '0', '1', "10", "110", "001", "000", '0', '-', "00"), -- i=1035
      ("1010100001100001", '1', '1', "10", "110", "001", "000", '0', '-', "00"), -- i=1036
      ("1010100001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1037
      ("1011000001100001", '0', '1', "11", "110", "001", "000", '0', '-', "00"), -- i=1038
      ("1011100001100001", '1', '1', "11", "110", "001", "000", '0', '-', "00"), -- i=1039
      ("1011100001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1040
      ("0101000001100000", '0', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1041
      ("0101100001100000", '1', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1042
      ("0101100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1043
      ("0100000001100000", '0', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1044
      ("0100100001100000", '1', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1045
      ("0100100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1046
      ("0000000010111001", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1047
      ("0000100010111001", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1048
      ("0000100010111001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1049
      ("1000000001100010", '0', '1', "00", "110", "010", "000", '0', '-', "00"), -- i=1050
      ("1000100001100010", '1', '1', "00", "110", "010", "000", '0', '-', "00"), -- i=1051
      ("1000100001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1052
      ("1001000001100010", '0', '1', "01", "110", "010", "000", '0', '-', "00"), -- i=1053
      ("1001100001100010", '1', '1', "01", "110", "010", "000", '0', '-', "00"), -- i=1054
      ("1001100001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1055
      ("1010000001100010", '0', '1', "10", "110", "010", "000", '0', '-', "00"), -- i=1056
      ("1010100001100010", '1', '1', "10", "110", "010", "000", '0', '-', "00"), -- i=1057
      ("1010100001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1058
      ("1011000001100010", '0', '1', "11", "110", "010", "000", '0', '-', "00"), -- i=1059
      ("1011100001100010", '1', '1', "11", "110", "010", "000", '0', '-', "00"), -- i=1060
      ("1011100001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1061
      ("0101000001100000", '0', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1062
      ("0101100001100000", '1', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1063
      ("0101100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1064
      ("0100000001100000", '0', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1065
      ("0100100001100000", '1', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1066
      ("0100100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1067
      ("0000000010000101", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1068
      ("0000100010000101", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1069
      ("0000100010000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1070
      ("1000000001100011", '0', '1', "00", "110", "011", "000", '0', '-', "00"), -- i=1071
      ("1000100001100011", '1', '1', "00", "110", "011", "000", '0', '-', "00"), -- i=1072
      ("1000100001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1073
      ("1001000001100011", '0', '1', "01", "110", "011", "000", '0', '-', "00"), -- i=1074
      ("1001100001100011", '1', '1', "01", "110", "011", "000", '0', '-', "00"), -- i=1075
      ("1001100001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1076
      ("1010000001100011", '0', '1', "10", "110", "011", "000", '0', '-', "00"), -- i=1077
      ("1010100001100011", '1', '1', "10", "110", "011", "000", '0', '-', "00"), -- i=1078
      ("1010100001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1079
      ("1011000001100011", '0', '1', "11", "110", "011", "000", '0', '-', "00"), -- i=1080
      ("1011100001100011", '1', '1', "11", "110", "011", "000", '0', '-', "00"), -- i=1081
      ("1011100001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1082
      ("0101000001100000", '0', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1083
      ("0101100001100000", '1', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1084
      ("0101100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1085
      ("0100000001100000", '0', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1086
      ("0100100001100000", '1', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1087
      ("0100100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1088
      ("0000000011100111", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1089
      ("0000100011100111", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1090
      ("0000100011100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1091
      ("1000000001100100", '0', '1', "00", "110", "100", "000", '0', '-', "00"), -- i=1092
      ("1000100001100100", '1', '1', "00", "110", "100", "000", '0', '-', "00"), -- i=1093
      ("1000100001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1094
      ("1001000001100100", '0', '1', "01", "110", "100", "000", '0', '-', "00"), -- i=1095
      ("1001100001100100", '1', '1', "01", "110", "100", "000", '0', '-', "00"), -- i=1096
      ("1001100001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1097
      ("1010000001100100", '0', '1', "10", "110", "100", "000", '0', '-', "00"), -- i=1098
      ("1010100001100100", '1', '1', "10", "110", "100", "000", '0', '-', "00"), -- i=1099
      ("1010100001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1100
      ("1011000001100100", '0', '1', "11", "110", "100", "000", '0', '-', "00"), -- i=1101
      ("1011100001100100", '1', '1', "11", "110", "100", "000", '0', '-', "00"), -- i=1102
      ("1011100001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1103
      ("0101000001100000", '0', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1104
      ("0101100001100000", '1', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1105
      ("0101100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1106
      ("0100000001100000", '0', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1107
      ("0100100001100000", '1', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1108
      ("0100100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1109
      ("0000000011011011", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1110
      ("0000100011011011", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1111
      ("0000100011011011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1112
      ("1000000001100101", '0', '1', "00", "110", "101", "000", '0', '-', "00"), -- i=1113
      ("1000100001100101", '1', '1', "00", "110", "101", "000", '0', '-', "00"), -- i=1114
      ("1000100001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1115
      ("1001000001100101", '0', '1', "01", "110", "101", "000", '0', '-', "00"), -- i=1116
      ("1001100001100101", '1', '1', "01", "110", "101", "000", '0', '-', "00"), -- i=1117
      ("1001100001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1118
      ("1010000001100101", '0', '1', "10", "110", "101", "000", '0', '-', "00"), -- i=1119
      ("1010100001100101", '1', '1', "10", "110", "101", "000", '0', '-', "00"), -- i=1120
      ("1010100001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1121
      ("1011000001100101", '0', '1', "11", "110", "101", "000", '0', '-', "00"), -- i=1122
      ("1011100001100101", '1', '1', "11", "110", "101", "000", '0', '-', "00"), -- i=1123
      ("1011100001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1124
      ("0101000001100000", '0', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1125
      ("0101100001100000", '1', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1126
      ("0101100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1127
      ("0100000001100000", '0', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1128
      ("0100100001100000", '1', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1129
      ("0100100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1130
      ("0000000000111100", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1131
      ("0000100000111100", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1132
      ("0000100000111100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1133
      ("1000000001100110", '0', '1', "00", "110", "110", "000", '0', '-', "00"), -- i=1134
      ("1000100001100110", '1', '1', "00", "110", "110", "000", '0', '-', "00"), -- i=1135
      ("1000100001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1136
      ("1001000001100110", '0', '1', "01", "110", "110", "000", '0', '-', "00"), -- i=1137
      ("1001100001100110", '1', '1', "01", "110", "110", "000", '0', '-', "00"), -- i=1138
      ("1001100001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1139
      ("1010000001100110", '0', '1', "10", "110", "110", "000", '0', '-', "00"), -- i=1140
      ("1010100001100110", '1', '1', "10", "110", "110", "000", '0', '-', "00"), -- i=1141
      ("1010100001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1142
      ("1011000001100110", '0', '1', "11", "110", "110", "000", '0', '-', "00"), -- i=1143
      ("1011100001100110", '1', '1', "11", "110", "110", "000", '0', '-', "00"), -- i=1144
      ("1011100001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1145
      ("0101000001100000", '0', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1146
      ("0101100001100000", '1', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1147
      ("0101100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1148
      ("0100000001100000", '0', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1149
      ("0100100001100000", '1', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1150
      ("0100100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1151
      ("0000000010111111", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1152
      ("0000100010111111", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1153
      ("0000100010111111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1154
      ("1000000001100111", '0', '1', "00", "110", "111", "000", '0', '-', "00"), -- i=1155
      ("1000100001100111", '1', '1', "00", "110", "111", "000", '0', '-', "00"), -- i=1156
      ("1000100001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1157
      ("1001000001100111", '0', '1', "01", "110", "111", "000", '0', '-', "00"), -- i=1158
      ("1001100001100111", '1', '1', "01", "110", "111", "000", '0', '-', "00"), -- i=1159
      ("1001100001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1160
      ("1010000001100111", '0', '1', "10", "110", "111", "000", '0', '-', "00"), -- i=1161
      ("1010100001100111", '1', '1', "10", "110", "111", "000", '0', '-', "00"), -- i=1162
      ("1010100001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1163
      ("1011000001100111", '0', '1', "11", "110", "111", "000", '0', '-', "00"), -- i=1164
      ("1011100001100111", '1', '1', "11", "110", "111", "000", '0', '-', "00"), -- i=1165
      ("1011100001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1166
      ("0101000001100000", '0', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1167
      ("0101100001100000", '1', '1', "--", "110", "---", "000", '0', '1', "01"), -- i=1168
      ("0101100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1169
      ("0100000001100000", '0', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1170
      ("0100100001100000", '1', '0', "--", "110", "000", "---", '1', '-', "--"), -- i=1171
      ("0100100001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1172
      ("0000000010001000", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1173
      ("0000100010001000", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1174
      ("0000100010001000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1175
      ("1000000001110000", '0', '1', "00", "111", "000", "000", '0', '-', "00"), -- i=1176
      ("1000100001110000", '1', '1', "00", "111", "000", "000", '0', '-', "00"), -- i=1177
      ("1000100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1178
      ("1001000001110000", '0', '1', "01", "111", "000", "000", '0', '-', "00"), -- i=1179
      ("1001100001110000", '1', '1', "01", "111", "000", "000", '0', '-', "00"), -- i=1180
      ("1001100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1181
      ("1010000001110000", '0', '1', "10", "111", "000", "000", '0', '-', "00"), -- i=1182
      ("1010100001110000", '1', '1', "10", "111", "000", "000", '0', '-', "00"), -- i=1183
      ("1010100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1184
      ("1011000001110000", '0', '1', "11", "111", "000", "000", '0', '-', "00"), -- i=1185
      ("1011100001110000", '1', '1', "11", "111", "000", "000", '0', '-', "00"), -- i=1186
      ("1011100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1187
      ("0101000001110000", '0', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1188
      ("0101100001110000", '1', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1189
      ("0101100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1190
      ("0100000001110000", '0', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1191
      ("0100100001110000", '1', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1192
      ("0100100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1193
      ("0000000000000011", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1194
      ("0000100000000011", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1195
      ("0000100000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1196
      ("1000000001110001", '0', '1', "00", "111", "001", "000", '0', '-', "00"), -- i=1197
      ("1000100001110001", '1', '1', "00", "111", "001", "000", '0', '-', "00"), -- i=1198
      ("1000100001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1199
      ("1001000001110001", '0', '1', "01", "111", "001", "000", '0', '-', "00"), -- i=1200
      ("1001100001110001", '1', '1', "01", "111", "001", "000", '0', '-', "00"), -- i=1201
      ("1001100001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1202
      ("1010000001110001", '0', '1', "10", "111", "001", "000", '0', '-', "00"), -- i=1203
      ("1010100001110001", '1', '1', "10", "111", "001", "000", '0', '-', "00"), -- i=1204
      ("1010100001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1205
      ("1011000001110001", '0', '1', "11", "111", "001", "000", '0', '-', "00"), -- i=1206
      ("1011100001110001", '1', '1', "11", "111", "001", "000", '0', '-', "00"), -- i=1207
      ("1011100001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1208
      ("0101000001110000", '0', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1209
      ("0101100001110000", '1', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1210
      ("0101100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1211
      ("0100000001110000", '0', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1212
      ("0100100001110000", '1', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1213
      ("0100100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1214
      ("0000000011111111", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1215
      ("0000100011111111", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1216
      ("0000100011111111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1217
      ("1000000001110010", '0', '1', "00", "111", "010", "000", '0', '-', "00"), -- i=1218
      ("1000100001110010", '1', '1', "00", "111", "010", "000", '0', '-', "00"), -- i=1219
      ("1000100001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1220
      ("1001000001110010", '0', '1', "01", "111", "010", "000", '0', '-', "00"), -- i=1221
      ("1001100001110010", '1', '1', "01", "111", "010", "000", '0', '-', "00"), -- i=1222
      ("1001100001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1223
      ("1010000001110010", '0', '1', "10", "111", "010", "000", '0', '-', "00"), -- i=1224
      ("1010100001110010", '1', '1', "10", "111", "010", "000", '0', '-', "00"), -- i=1225
      ("1010100001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1226
      ("1011000001110010", '0', '1', "11", "111", "010", "000", '0', '-', "00"), -- i=1227
      ("1011100001110010", '1', '1', "11", "111", "010", "000", '0', '-', "00"), -- i=1228
      ("1011100001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1229
      ("0101000001110000", '0', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1230
      ("0101100001110000", '1', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1231
      ("0101100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1232
      ("0100000001110000", '0', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1233
      ("0100100001110000", '1', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1234
      ("0100100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1235
      ("0000000001011010", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1236
      ("0000100001011010", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1237
      ("0000100001011010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1238
      ("1000000001110011", '0', '1', "00", "111", "011", "000", '0', '-', "00"), -- i=1239
      ("1000100001110011", '1', '1', "00", "111", "011", "000", '0', '-', "00"), -- i=1240
      ("1000100001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1241
      ("1001000001110011", '0', '1', "01", "111", "011", "000", '0', '-', "00"), -- i=1242
      ("1001100001110011", '1', '1', "01", "111", "011", "000", '0', '-', "00"), -- i=1243
      ("1001100001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1244
      ("1010000001110011", '0', '1', "10", "111", "011", "000", '0', '-', "00"), -- i=1245
      ("1010100001110011", '1', '1', "10", "111", "011", "000", '0', '-', "00"), -- i=1246
      ("1010100001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1247
      ("1011000001110011", '0', '1', "11", "111", "011", "000", '0', '-', "00"), -- i=1248
      ("1011100001110011", '1', '1', "11", "111", "011", "000", '0', '-', "00"), -- i=1249
      ("1011100001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1250
      ("0101000001110000", '0', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1251
      ("0101100001110000", '1', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1252
      ("0101100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1253
      ("0100000001110000", '0', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1254
      ("0100100001110000", '1', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1255
      ("0100100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1256
      ("0000000010010000", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1257
      ("0000100010010000", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1258
      ("0000100010010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1259
      ("1000000001110100", '0', '1', "00", "111", "100", "000", '0', '-', "00"), -- i=1260
      ("1000100001110100", '1', '1', "00", "111", "100", "000", '0', '-', "00"), -- i=1261
      ("1000100001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1262
      ("1001000001110100", '0', '1', "01", "111", "100", "000", '0', '-', "00"), -- i=1263
      ("1001100001110100", '1', '1', "01", "111", "100", "000", '0', '-', "00"), -- i=1264
      ("1001100001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1265
      ("1010000001110100", '0', '1', "10", "111", "100", "000", '0', '-', "00"), -- i=1266
      ("1010100001110100", '1', '1', "10", "111", "100", "000", '0', '-', "00"), -- i=1267
      ("1010100001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1268
      ("1011000001110100", '0', '1', "11", "111", "100", "000", '0', '-', "00"), -- i=1269
      ("1011100001110100", '1', '1', "11", "111", "100", "000", '0', '-', "00"), -- i=1270
      ("1011100001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1271
      ("0101000001110000", '0', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1272
      ("0101100001110000", '1', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1273
      ("0101100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1274
      ("0100000001110000", '0', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1275
      ("0100100001110000", '1', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1276
      ("0100100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1277
      ("0000000001111010", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1278
      ("0000100001111010", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1279
      ("0000100001111010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1280
      ("1000000001110101", '0', '1', "00", "111", "101", "000", '0', '-', "00"), -- i=1281
      ("1000100001110101", '1', '1', "00", "111", "101", "000", '0', '-', "00"), -- i=1282
      ("1000100001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1283
      ("1001000001110101", '0', '1', "01", "111", "101", "000", '0', '-', "00"), -- i=1284
      ("1001100001110101", '1', '1', "01", "111", "101", "000", '0', '-', "00"), -- i=1285
      ("1001100001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1286
      ("1010000001110101", '0', '1', "10", "111", "101", "000", '0', '-', "00"), -- i=1287
      ("1010100001110101", '1', '1', "10", "111", "101", "000", '0', '-', "00"), -- i=1288
      ("1010100001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1289
      ("1011000001110101", '0', '1', "11", "111", "101", "000", '0', '-', "00"), -- i=1290
      ("1011100001110101", '1', '1', "11", "111", "101", "000", '0', '-', "00"), -- i=1291
      ("1011100001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1292
      ("0101000001110000", '0', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1293
      ("0101100001110000", '1', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1294
      ("0101100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1295
      ("0100000001110000", '0', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1296
      ("0100100001110000", '1', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1297
      ("0100100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1298
      ("0000000011000100", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1299
      ("0000100011000100", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1300
      ("0000100011000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1301
      ("1000000001110110", '0', '1', "00", "111", "110", "000", '0', '-', "00"), -- i=1302
      ("1000100001110110", '1', '1', "00", "111", "110", "000", '0', '-', "00"), -- i=1303
      ("1000100001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1304
      ("1001000001110110", '0', '1', "01", "111", "110", "000", '0', '-', "00"), -- i=1305
      ("1001100001110110", '1', '1', "01", "111", "110", "000", '0', '-', "00"), -- i=1306
      ("1001100001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1307
      ("1010000001110110", '0', '1', "10", "111", "110", "000", '0', '-', "00"), -- i=1308
      ("1010100001110110", '1', '1', "10", "111", "110", "000", '0', '-', "00"), -- i=1309
      ("1010100001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1310
      ("1011000001110110", '0', '1', "11", "111", "110", "000", '0', '-', "00"), -- i=1311
      ("1011100001110110", '1', '1', "11", "111", "110", "000", '0', '-', "00"), -- i=1312
      ("1011100001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1313
      ("0101000001110000", '0', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1314
      ("0101100001110000", '1', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1315
      ("0101100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1316
      ("0100000001110000", '0', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1317
      ("0100100001110000", '1', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1318
      ("0100100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1319
      ("0000000010101000", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1320
      ("0000100010101000", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1321
      ("0000100010101000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1322
      ("1000000001110111", '0', '1', "00", "111", "111", "000", '0', '-', "00"), -- i=1323
      ("1000100001110111", '1', '1', "00", "111", "111", "000", '0', '-', "00"), -- i=1324
      ("1000100001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1325
      ("1001000001110111", '0', '1', "01", "111", "111", "000", '0', '-', "00"), -- i=1326
      ("1001100001110111", '1', '1', "01", "111", "111", "000", '0', '-', "00"), -- i=1327
      ("1001100001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1328
      ("1010000001110111", '0', '1', "10", "111", "111", "000", '0', '-', "00"), -- i=1329
      ("1010100001110111", '1', '1', "10", "111", "111", "000", '0', '-', "00"), -- i=1330
      ("1010100001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1331
      ("1011000001110111", '0', '1', "11", "111", "111", "000", '0', '-', "00"), -- i=1332
      ("1011100001110111", '1', '1', "11", "111", "111", "000", '0', '-', "00"), -- i=1333
      ("1011100001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1334
      ("0101000001110000", '0', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1335
      ("0101100001110000", '1', '1', "--", "111", "---", "000", '0', '1', "01"), -- i=1336
      ("0101100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1337
      ("0100000001110000", '0', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1338
      ("0100100001110000", '1', '0', "--", "111", "000", "---", '1', '-', "--"), -- i=1339
      ("0100100001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1340
      ("0000000001100010", '0', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1341
      ("0000100001100010", '1', '1', "--", "---", "---", "000", '0', '-', "10"), -- i=1342
      ("0000100001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1343
      ("1000000100000000", '0', '1', "00", "000", "000", "001", '0', '-', "00"), -- i=1344
      ("1000100100000000", '1', '1', "00", "000", "000", "001", '0', '-', "00"), -- i=1345
      ("1000100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1346
      ("1001000100000000", '0', '1', "01", "000", "000", "001", '0', '-', "00"), -- i=1347
      ("1001100100000000", '1', '1', "01", "000", "000", "001", '0', '-', "00"), -- i=1348
      ("1001100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1349
      ("1010000100000000", '0', '1', "10", "000", "000", "001", '0', '-', "00"), -- i=1350
      ("1010100100000000", '1', '1', "10", "000", "000", "001", '0', '-', "00"), -- i=1351
      ("1010100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1352
      ("1011000100000000", '0', '1', "11", "000", "000", "001", '0', '-', "00"), -- i=1353
      ("1011100100000000", '1', '1', "11", "000", "000", "001", '0', '-', "00"), -- i=1354
      ("1011100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1355
      ("0101000100000000", '0', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1356
      ("0101100100000000", '1', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1357
      ("0101100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1358
      ("0100000100000000", '0', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1359
      ("0100100100000000", '1', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1360
      ("0100100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1361
      ("0000000110011100", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1362
      ("0000100110011100", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1363
      ("0000100110011100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1364
      ("1000000100000001", '0', '1', "00", "000", "001", "001", '0', '-', "00"), -- i=1365
      ("1000100100000001", '1', '1', "00", "000", "001", "001", '0', '-', "00"), -- i=1366
      ("1000100100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1367
      ("1001000100000001", '0', '1', "01", "000", "001", "001", '0', '-', "00"), -- i=1368
      ("1001100100000001", '1', '1', "01", "000", "001", "001", '0', '-', "00"), -- i=1369
      ("1001100100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1370
      ("1010000100000001", '0', '1', "10", "000", "001", "001", '0', '-', "00"), -- i=1371
      ("1010100100000001", '1', '1', "10", "000", "001", "001", '0', '-', "00"), -- i=1372
      ("1010100100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1373
      ("1011000100000001", '0', '1', "11", "000", "001", "001", '0', '-', "00"), -- i=1374
      ("1011100100000001", '1', '1', "11", "000", "001", "001", '0', '-', "00"), -- i=1375
      ("1011100100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1376
      ("0101000100000000", '0', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1377
      ("0101100100000000", '1', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1378
      ("0101100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1379
      ("0100000100000000", '0', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1380
      ("0100100100000000", '1', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1381
      ("0100100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1382
      ("0000000101111111", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1383
      ("0000100101111111", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1384
      ("0000100101111111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1385
      ("1000000100000010", '0', '1', "00", "000", "010", "001", '0', '-', "00"), -- i=1386
      ("1000100100000010", '1', '1', "00", "000", "010", "001", '0', '-', "00"), -- i=1387
      ("1000100100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1388
      ("1001000100000010", '0', '1', "01", "000", "010", "001", '0', '-', "00"), -- i=1389
      ("1001100100000010", '1', '1', "01", "000", "010", "001", '0', '-', "00"), -- i=1390
      ("1001100100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1391
      ("1010000100000010", '0', '1', "10", "000", "010", "001", '0', '-', "00"), -- i=1392
      ("1010100100000010", '1', '1', "10", "000", "010", "001", '0', '-', "00"), -- i=1393
      ("1010100100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1394
      ("1011000100000010", '0', '1', "11", "000", "010", "001", '0', '-', "00"), -- i=1395
      ("1011100100000010", '1', '1', "11", "000", "010", "001", '0', '-', "00"), -- i=1396
      ("1011100100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1397
      ("0101000100000000", '0', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1398
      ("0101100100000000", '1', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1399
      ("0101100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1400
      ("0100000100000000", '0', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1401
      ("0100100100000000", '1', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1402
      ("0100100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1403
      ("0000000100110111", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1404
      ("0000100100110111", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1405
      ("0000100100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1406
      ("1000000100000011", '0', '1', "00", "000", "011", "001", '0', '-', "00"), -- i=1407
      ("1000100100000011", '1', '1', "00", "000", "011", "001", '0', '-', "00"), -- i=1408
      ("1000100100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1409
      ("1001000100000011", '0', '1', "01", "000", "011", "001", '0', '-', "00"), -- i=1410
      ("1001100100000011", '1', '1', "01", "000", "011", "001", '0', '-', "00"), -- i=1411
      ("1001100100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1412
      ("1010000100000011", '0', '1', "10", "000", "011", "001", '0', '-', "00"), -- i=1413
      ("1010100100000011", '1', '1', "10", "000", "011", "001", '0', '-', "00"), -- i=1414
      ("1010100100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1415
      ("1011000100000011", '0', '1', "11", "000", "011", "001", '0', '-', "00"), -- i=1416
      ("1011100100000011", '1', '1', "11", "000", "011", "001", '0', '-', "00"), -- i=1417
      ("1011100100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1418
      ("0101000100000000", '0', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1419
      ("0101100100000000", '1', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1420
      ("0101100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1421
      ("0100000100000000", '0', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1422
      ("0100100100000000", '1', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1423
      ("0100100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1424
      ("0000000101101100", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1425
      ("0000100101101100", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1426
      ("0000100101101100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1427
      ("1000000100000100", '0', '1', "00", "000", "100", "001", '0', '-', "00"), -- i=1428
      ("1000100100000100", '1', '1', "00", "000", "100", "001", '0', '-', "00"), -- i=1429
      ("1000100100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1430
      ("1001000100000100", '0', '1', "01", "000", "100", "001", '0', '-', "00"), -- i=1431
      ("1001100100000100", '1', '1', "01", "000", "100", "001", '0', '-', "00"), -- i=1432
      ("1001100100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1433
      ("1010000100000100", '0', '1', "10", "000", "100", "001", '0', '-', "00"), -- i=1434
      ("1010100100000100", '1', '1', "10", "000", "100", "001", '0', '-', "00"), -- i=1435
      ("1010100100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1436
      ("1011000100000100", '0', '1', "11", "000", "100", "001", '0', '-', "00"), -- i=1437
      ("1011100100000100", '1', '1', "11", "000", "100", "001", '0', '-', "00"), -- i=1438
      ("1011100100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1439
      ("0101000100000000", '0', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1440
      ("0101100100000000", '1', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1441
      ("0101100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1442
      ("0100000100000000", '0', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1443
      ("0100100100000000", '1', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1444
      ("0100100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1445
      ("0000000100011011", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1446
      ("0000100100011011", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1447
      ("0000100100011011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1448
      ("1000000100000101", '0', '1', "00", "000", "101", "001", '0', '-', "00"), -- i=1449
      ("1000100100000101", '1', '1', "00", "000", "101", "001", '0', '-', "00"), -- i=1450
      ("1000100100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1451
      ("1001000100000101", '0', '1', "01", "000", "101", "001", '0', '-', "00"), -- i=1452
      ("1001100100000101", '1', '1', "01", "000", "101", "001", '0', '-', "00"), -- i=1453
      ("1001100100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1454
      ("1010000100000101", '0', '1', "10", "000", "101", "001", '0', '-', "00"), -- i=1455
      ("1010100100000101", '1', '1', "10", "000", "101", "001", '0', '-', "00"), -- i=1456
      ("1010100100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1457
      ("1011000100000101", '0', '1', "11", "000", "101", "001", '0', '-', "00"), -- i=1458
      ("1011100100000101", '1', '1', "11", "000", "101", "001", '0', '-', "00"), -- i=1459
      ("1011100100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1460
      ("0101000100000000", '0', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1461
      ("0101100100000000", '1', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1462
      ("0101100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1463
      ("0100000100000000", '0', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1464
      ("0100100100000000", '1', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1465
      ("0100100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1466
      ("0000000110001111", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1467
      ("0000100110001111", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1468
      ("0000100110001111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1469
      ("1000000100000110", '0', '1', "00", "000", "110", "001", '0', '-', "00"), -- i=1470
      ("1000100100000110", '1', '1', "00", "000", "110", "001", '0', '-', "00"), -- i=1471
      ("1000100100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1472
      ("1001000100000110", '0', '1', "01", "000", "110", "001", '0', '-', "00"), -- i=1473
      ("1001100100000110", '1', '1', "01", "000", "110", "001", '0', '-', "00"), -- i=1474
      ("1001100100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1475
      ("1010000100000110", '0', '1', "10", "000", "110", "001", '0', '-', "00"), -- i=1476
      ("1010100100000110", '1', '1', "10", "000", "110", "001", '0', '-', "00"), -- i=1477
      ("1010100100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1478
      ("1011000100000110", '0', '1', "11", "000", "110", "001", '0', '-', "00"), -- i=1479
      ("1011100100000110", '1', '1', "11", "000", "110", "001", '0', '-', "00"), -- i=1480
      ("1011100100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1481
      ("0101000100000000", '0', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1482
      ("0101100100000000", '1', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1483
      ("0101100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1484
      ("0100000100000000", '0', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1485
      ("0100100100000000", '1', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1486
      ("0100100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1487
      ("0000000101100000", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1488
      ("0000100101100000", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1489
      ("0000100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1490
      ("1000000100000111", '0', '1', "00", "000", "111", "001", '0', '-', "00"), -- i=1491
      ("1000100100000111", '1', '1', "00", "000", "111", "001", '0', '-', "00"), -- i=1492
      ("1000100100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1493
      ("1001000100000111", '0', '1', "01", "000", "111", "001", '0', '-', "00"), -- i=1494
      ("1001100100000111", '1', '1', "01", "000", "111", "001", '0', '-', "00"), -- i=1495
      ("1001100100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1496
      ("1010000100000111", '0', '1', "10", "000", "111", "001", '0', '-', "00"), -- i=1497
      ("1010100100000111", '1', '1', "10", "000", "111", "001", '0', '-', "00"), -- i=1498
      ("1010100100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1499
      ("1011000100000111", '0', '1', "11", "000", "111", "001", '0', '-', "00"), -- i=1500
      ("1011100100000111", '1', '1', "11", "000", "111", "001", '0', '-', "00"), -- i=1501
      ("1011100100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1502
      ("0101000100000000", '0', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1503
      ("0101100100000000", '1', '1', "--", "000", "---", "001", '0', '1', "01"), -- i=1504
      ("0101100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1505
      ("0100000100000000", '0', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1506
      ("0100100100000000", '1', '0', "--", "000", "001", "---", '1', '-', "--"), -- i=1507
      ("0100100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1508
      ("0000000101111111", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1509
      ("0000100101111111", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1510
      ("0000100101111111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1511
      ("1000000100010000", '0', '1', "00", "001", "000", "001", '0', '-', "00"), -- i=1512
      ("1000100100010000", '1', '1', "00", "001", "000", "001", '0', '-', "00"), -- i=1513
      ("1000100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1514
      ("1001000100010000", '0', '1', "01", "001", "000", "001", '0', '-', "00"), -- i=1515
      ("1001100100010000", '1', '1', "01", "001", "000", "001", '0', '-', "00"), -- i=1516
      ("1001100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1517
      ("1010000100010000", '0', '1', "10", "001", "000", "001", '0', '-', "00"), -- i=1518
      ("1010100100010000", '1', '1', "10", "001", "000", "001", '0', '-', "00"), -- i=1519
      ("1010100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1520
      ("1011000100010000", '0', '1', "11", "001", "000", "001", '0', '-', "00"), -- i=1521
      ("1011100100010000", '1', '1', "11", "001", "000", "001", '0', '-', "00"), -- i=1522
      ("1011100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1523
      ("0101000100010000", '0', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1524
      ("0101100100010000", '1', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1525
      ("0101100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1526
      ("0100000100010000", '0', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1527
      ("0100100100010000", '1', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1528
      ("0100100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1529
      ("0000000100101111", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1530
      ("0000100100101111", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1531
      ("0000100100101111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1532
      ("1000000100010001", '0', '1', "00", "001", "001", "001", '0', '-', "00"), -- i=1533
      ("1000100100010001", '1', '1', "00", "001", "001", "001", '0', '-', "00"), -- i=1534
      ("1000100100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1535
      ("1001000100010001", '0', '1', "01", "001", "001", "001", '0', '-', "00"), -- i=1536
      ("1001100100010001", '1', '1', "01", "001", "001", "001", '0', '-', "00"), -- i=1537
      ("1001100100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1538
      ("1010000100010001", '0', '1', "10", "001", "001", "001", '0', '-', "00"), -- i=1539
      ("1010100100010001", '1', '1', "10", "001", "001", "001", '0', '-', "00"), -- i=1540
      ("1010100100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1541
      ("1011000100010001", '0', '1', "11", "001", "001", "001", '0', '-', "00"), -- i=1542
      ("1011100100010001", '1', '1', "11", "001", "001", "001", '0', '-', "00"), -- i=1543
      ("1011100100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1544
      ("0101000100010000", '0', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1545
      ("0101100100010000", '1', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1546
      ("0101100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1547
      ("0100000100010000", '0', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1548
      ("0100100100010000", '1', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1549
      ("0100100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1550
      ("0000000100100101", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1551
      ("0000100100100101", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1552
      ("0000100100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1553
      ("1000000100010010", '0', '1', "00", "001", "010", "001", '0', '-', "00"), -- i=1554
      ("1000100100010010", '1', '1', "00", "001", "010", "001", '0', '-', "00"), -- i=1555
      ("1000100100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1556
      ("1001000100010010", '0', '1', "01", "001", "010", "001", '0', '-', "00"), -- i=1557
      ("1001100100010010", '1', '1', "01", "001", "010", "001", '0', '-', "00"), -- i=1558
      ("1001100100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1559
      ("1010000100010010", '0', '1', "10", "001", "010", "001", '0', '-', "00"), -- i=1560
      ("1010100100010010", '1', '1', "10", "001", "010", "001", '0', '-', "00"), -- i=1561
      ("1010100100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1562
      ("1011000100010010", '0', '1', "11", "001", "010", "001", '0', '-', "00"), -- i=1563
      ("1011100100010010", '1', '1', "11", "001", "010", "001", '0', '-', "00"), -- i=1564
      ("1011100100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1565
      ("0101000100010000", '0', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1566
      ("0101100100010000", '1', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1567
      ("0101100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1568
      ("0100000100010000", '0', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1569
      ("0100100100010000", '1', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1570
      ("0100100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1571
      ("0000000101000010", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1572
      ("0000100101000010", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1573
      ("0000100101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1574
      ("1000000100010011", '0', '1', "00", "001", "011", "001", '0', '-', "00"), -- i=1575
      ("1000100100010011", '1', '1', "00", "001", "011", "001", '0', '-', "00"), -- i=1576
      ("1000100100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1577
      ("1001000100010011", '0', '1', "01", "001", "011", "001", '0', '-', "00"), -- i=1578
      ("1001100100010011", '1', '1', "01", "001", "011", "001", '0', '-', "00"), -- i=1579
      ("1001100100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1580
      ("1010000100010011", '0', '1', "10", "001", "011", "001", '0', '-', "00"), -- i=1581
      ("1010100100010011", '1', '1', "10", "001", "011", "001", '0', '-', "00"), -- i=1582
      ("1010100100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1583
      ("1011000100010011", '0', '1', "11", "001", "011", "001", '0', '-', "00"), -- i=1584
      ("1011100100010011", '1', '1', "11", "001", "011", "001", '0', '-', "00"), -- i=1585
      ("1011100100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1586
      ("0101000100010000", '0', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1587
      ("0101100100010000", '1', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1588
      ("0101100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1589
      ("0100000100010000", '0', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1590
      ("0100100100010000", '1', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1591
      ("0100100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1592
      ("0000000101111110", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1593
      ("0000100101111110", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1594
      ("0000100101111110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1595
      ("1000000100010100", '0', '1', "00", "001", "100", "001", '0', '-', "00"), -- i=1596
      ("1000100100010100", '1', '1', "00", "001", "100", "001", '0', '-', "00"), -- i=1597
      ("1000100100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1598
      ("1001000100010100", '0', '1', "01", "001", "100", "001", '0', '-', "00"), -- i=1599
      ("1001100100010100", '1', '1', "01", "001", "100", "001", '0', '-', "00"), -- i=1600
      ("1001100100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1601
      ("1010000100010100", '0', '1', "10", "001", "100", "001", '0', '-', "00"), -- i=1602
      ("1010100100010100", '1', '1', "10", "001", "100", "001", '0', '-', "00"), -- i=1603
      ("1010100100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1604
      ("1011000100010100", '0', '1', "11", "001", "100", "001", '0', '-', "00"), -- i=1605
      ("1011100100010100", '1', '1', "11", "001", "100", "001", '0', '-', "00"), -- i=1606
      ("1011100100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1607
      ("0101000100010000", '0', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1608
      ("0101100100010000", '1', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1609
      ("0101100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1610
      ("0100000100010000", '0', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1611
      ("0100100100010000", '1', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1612
      ("0100100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1613
      ("0000000101010110", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1614
      ("0000100101010110", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1615
      ("0000100101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1616
      ("1000000100010101", '0', '1', "00", "001", "101", "001", '0', '-', "00"), -- i=1617
      ("1000100100010101", '1', '1', "00", "001", "101", "001", '0', '-', "00"), -- i=1618
      ("1000100100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1619
      ("1001000100010101", '0', '1', "01", "001", "101", "001", '0', '-', "00"), -- i=1620
      ("1001100100010101", '1', '1', "01", "001", "101", "001", '0', '-', "00"), -- i=1621
      ("1001100100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1622
      ("1010000100010101", '0', '1', "10", "001", "101", "001", '0', '-', "00"), -- i=1623
      ("1010100100010101", '1', '1', "10", "001", "101", "001", '0', '-', "00"), -- i=1624
      ("1010100100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1625
      ("1011000100010101", '0', '1', "11", "001", "101", "001", '0', '-', "00"), -- i=1626
      ("1011100100010101", '1', '1', "11", "001", "101", "001", '0', '-', "00"), -- i=1627
      ("1011100100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1628
      ("0101000100010000", '0', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1629
      ("0101100100010000", '1', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1630
      ("0101100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1631
      ("0100000100010000", '0', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1632
      ("0100100100010000", '1', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1633
      ("0100100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1634
      ("0000000111111000", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1635
      ("0000100111111000", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1636
      ("0000100111111000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1637
      ("1000000100010110", '0', '1', "00", "001", "110", "001", '0', '-', "00"), -- i=1638
      ("1000100100010110", '1', '1', "00", "001", "110", "001", '0', '-', "00"), -- i=1639
      ("1000100100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1640
      ("1001000100010110", '0', '1', "01", "001", "110", "001", '0', '-', "00"), -- i=1641
      ("1001100100010110", '1', '1', "01", "001", "110", "001", '0', '-', "00"), -- i=1642
      ("1001100100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1643
      ("1010000100010110", '0', '1', "10", "001", "110", "001", '0', '-', "00"), -- i=1644
      ("1010100100010110", '1', '1', "10", "001", "110", "001", '0', '-', "00"), -- i=1645
      ("1010100100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1646
      ("1011000100010110", '0', '1', "11", "001", "110", "001", '0', '-', "00"), -- i=1647
      ("1011100100010110", '1', '1', "11", "001", "110", "001", '0', '-', "00"), -- i=1648
      ("1011100100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1649
      ("0101000100010000", '0', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1650
      ("0101100100010000", '1', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1651
      ("0101100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1652
      ("0100000100010000", '0', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1653
      ("0100100100010000", '1', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1654
      ("0100100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1655
      ("0000000100000110", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1656
      ("0000100100000110", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1657
      ("0000100100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1658
      ("1000000100010111", '0', '1', "00", "001", "111", "001", '0', '-', "00"), -- i=1659
      ("1000100100010111", '1', '1', "00", "001", "111", "001", '0', '-', "00"), -- i=1660
      ("1000100100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1661
      ("1001000100010111", '0', '1', "01", "001", "111", "001", '0', '-', "00"), -- i=1662
      ("1001100100010111", '1', '1', "01", "001", "111", "001", '0', '-', "00"), -- i=1663
      ("1001100100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1664
      ("1010000100010111", '0', '1', "10", "001", "111", "001", '0', '-', "00"), -- i=1665
      ("1010100100010111", '1', '1', "10", "001", "111", "001", '0', '-', "00"), -- i=1666
      ("1010100100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1667
      ("1011000100010111", '0', '1', "11", "001", "111", "001", '0', '-', "00"), -- i=1668
      ("1011100100010111", '1', '1', "11", "001", "111", "001", '0', '-', "00"), -- i=1669
      ("1011100100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1670
      ("0101000100010000", '0', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1671
      ("0101100100010000", '1', '1', "--", "001", "---", "001", '0', '1', "01"), -- i=1672
      ("0101100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1673
      ("0100000100010000", '0', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1674
      ("0100100100010000", '1', '0', "--", "001", "001", "---", '1', '-', "--"), -- i=1675
      ("0100100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1676
      ("0000000111100001", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1677
      ("0000100111100001", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1678
      ("0000100111100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1679
      ("1000000100100000", '0', '1', "00", "010", "000", "001", '0', '-', "00"), -- i=1680
      ("1000100100100000", '1', '1', "00", "010", "000", "001", '0', '-', "00"), -- i=1681
      ("1000100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1682
      ("1001000100100000", '0', '1', "01", "010", "000", "001", '0', '-', "00"), -- i=1683
      ("1001100100100000", '1', '1', "01", "010", "000", "001", '0', '-', "00"), -- i=1684
      ("1001100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1685
      ("1010000100100000", '0', '1', "10", "010", "000", "001", '0', '-', "00"), -- i=1686
      ("1010100100100000", '1', '1', "10", "010", "000", "001", '0', '-', "00"), -- i=1687
      ("1010100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1688
      ("1011000100100000", '0', '1', "11", "010", "000", "001", '0', '-', "00"), -- i=1689
      ("1011100100100000", '1', '1', "11", "010", "000", "001", '0', '-', "00"), -- i=1690
      ("1011100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1691
      ("0101000100100000", '0', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1692
      ("0101100100100000", '1', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1693
      ("0101100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1694
      ("0100000100100000", '0', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1695
      ("0100100100100000", '1', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1696
      ("0100100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1697
      ("0000000111001110", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1698
      ("0000100111001110", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1699
      ("0000100111001110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1700
      ("1000000100100001", '0', '1', "00", "010", "001", "001", '0', '-', "00"), -- i=1701
      ("1000100100100001", '1', '1', "00", "010", "001", "001", '0', '-', "00"), -- i=1702
      ("1000100100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1703
      ("1001000100100001", '0', '1', "01", "010", "001", "001", '0', '-', "00"), -- i=1704
      ("1001100100100001", '1', '1', "01", "010", "001", "001", '0', '-', "00"), -- i=1705
      ("1001100100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1706
      ("1010000100100001", '0', '1', "10", "010", "001", "001", '0', '-', "00"), -- i=1707
      ("1010100100100001", '1', '1', "10", "010", "001", "001", '0', '-', "00"), -- i=1708
      ("1010100100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1709
      ("1011000100100001", '0', '1', "11", "010", "001", "001", '0', '-', "00"), -- i=1710
      ("1011100100100001", '1', '1', "11", "010", "001", "001", '0', '-', "00"), -- i=1711
      ("1011100100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1712
      ("0101000100100000", '0', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1713
      ("0101100100100000", '1', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1714
      ("0101100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1715
      ("0100000100100000", '0', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1716
      ("0100100100100000", '1', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1717
      ("0100100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1718
      ("0000000110000111", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1719
      ("0000100110000111", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1720
      ("0000100110000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1721
      ("1000000100100010", '0', '1', "00", "010", "010", "001", '0', '-', "00"), -- i=1722
      ("1000100100100010", '1', '1', "00", "010", "010", "001", '0', '-', "00"), -- i=1723
      ("1000100100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1724
      ("1001000100100010", '0', '1', "01", "010", "010", "001", '0', '-', "00"), -- i=1725
      ("1001100100100010", '1', '1', "01", "010", "010", "001", '0', '-', "00"), -- i=1726
      ("1001100100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1727
      ("1010000100100010", '0', '1', "10", "010", "010", "001", '0', '-', "00"), -- i=1728
      ("1010100100100010", '1', '1', "10", "010", "010", "001", '0', '-', "00"), -- i=1729
      ("1010100100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1730
      ("1011000100100010", '0', '1', "11", "010", "010", "001", '0', '-', "00"), -- i=1731
      ("1011100100100010", '1', '1', "11", "010", "010", "001", '0', '-', "00"), -- i=1732
      ("1011100100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1733
      ("0101000100100000", '0', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1734
      ("0101100100100000", '1', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1735
      ("0101100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1736
      ("0100000100100000", '0', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1737
      ("0100100100100000", '1', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1738
      ("0100100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1739
      ("0000000100001000", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1740
      ("0000100100001000", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1741
      ("0000100100001000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1742
      ("1000000100100011", '0', '1', "00", "010", "011", "001", '0', '-', "00"), -- i=1743
      ("1000100100100011", '1', '1', "00", "010", "011", "001", '0', '-', "00"), -- i=1744
      ("1000100100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1745
      ("1001000100100011", '0', '1', "01", "010", "011", "001", '0', '-', "00"), -- i=1746
      ("1001100100100011", '1', '1', "01", "010", "011", "001", '0', '-', "00"), -- i=1747
      ("1001100100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1748
      ("1010000100100011", '0', '1', "10", "010", "011", "001", '0', '-', "00"), -- i=1749
      ("1010100100100011", '1', '1', "10", "010", "011", "001", '0', '-', "00"), -- i=1750
      ("1010100100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1751
      ("1011000100100011", '0', '1', "11", "010", "011", "001", '0', '-', "00"), -- i=1752
      ("1011100100100011", '1', '1', "11", "010", "011", "001", '0', '-', "00"), -- i=1753
      ("1011100100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1754
      ("0101000100100000", '0', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1755
      ("0101100100100000", '1', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1756
      ("0101100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1757
      ("0100000100100000", '0', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1758
      ("0100100100100000", '1', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1759
      ("0100100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1760
      ("0000000110011010", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1761
      ("0000100110011010", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1762
      ("0000100110011010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1763
      ("1000000100100100", '0', '1', "00", "010", "100", "001", '0', '-', "00"), -- i=1764
      ("1000100100100100", '1', '1', "00", "010", "100", "001", '0', '-', "00"), -- i=1765
      ("1000100100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1766
      ("1001000100100100", '0', '1', "01", "010", "100", "001", '0', '-', "00"), -- i=1767
      ("1001100100100100", '1', '1', "01", "010", "100", "001", '0', '-', "00"), -- i=1768
      ("1001100100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1769
      ("1010000100100100", '0', '1', "10", "010", "100", "001", '0', '-', "00"), -- i=1770
      ("1010100100100100", '1', '1', "10", "010", "100", "001", '0', '-', "00"), -- i=1771
      ("1010100100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1772
      ("1011000100100100", '0', '1', "11", "010", "100", "001", '0', '-', "00"), -- i=1773
      ("1011100100100100", '1', '1', "11", "010", "100", "001", '0', '-', "00"), -- i=1774
      ("1011100100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1775
      ("0101000100100000", '0', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1776
      ("0101100100100000", '1', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1777
      ("0101100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1778
      ("0100000100100000", '0', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1779
      ("0100100100100000", '1', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1780
      ("0100100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1781
      ("0000000111100000", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1782
      ("0000100111100000", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1783
      ("0000100111100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1784
      ("1000000100100101", '0', '1', "00", "010", "101", "001", '0', '-', "00"), -- i=1785
      ("1000100100100101", '1', '1', "00", "010", "101", "001", '0', '-', "00"), -- i=1786
      ("1000100100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1787
      ("1001000100100101", '0', '1', "01", "010", "101", "001", '0', '-', "00"), -- i=1788
      ("1001100100100101", '1', '1', "01", "010", "101", "001", '0', '-', "00"), -- i=1789
      ("1001100100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1790
      ("1010000100100101", '0', '1', "10", "010", "101", "001", '0', '-', "00"), -- i=1791
      ("1010100100100101", '1', '1', "10", "010", "101", "001", '0', '-', "00"), -- i=1792
      ("1010100100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1793
      ("1011000100100101", '0', '1', "11", "010", "101", "001", '0', '-', "00"), -- i=1794
      ("1011100100100101", '1', '1', "11", "010", "101", "001", '0', '-', "00"), -- i=1795
      ("1011100100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1796
      ("0101000100100000", '0', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1797
      ("0101100100100000", '1', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1798
      ("0101100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1799
      ("0100000100100000", '0', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1800
      ("0100100100100000", '1', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1801
      ("0100100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1802
      ("0000000100010000", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1803
      ("0000100100010000", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1804
      ("0000100100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1805
      ("1000000100100110", '0', '1', "00", "010", "110", "001", '0', '-', "00"), -- i=1806
      ("1000100100100110", '1', '1', "00", "010", "110", "001", '0', '-', "00"), -- i=1807
      ("1000100100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1808
      ("1001000100100110", '0', '1', "01", "010", "110", "001", '0', '-', "00"), -- i=1809
      ("1001100100100110", '1', '1', "01", "010", "110", "001", '0', '-', "00"), -- i=1810
      ("1001100100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1811
      ("1010000100100110", '0', '1', "10", "010", "110", "001", '0', '-', "00"), -- i=1812
      ("1010100100100110", '1', '1', "10", "010", "110", "001", '0', '-', "00"), -- i=1813
      ("1010100100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1814
      ("1011000100100110", '0', '1', "11", "010", "110", "001", '0', '-', "00"), -- i=1815
      ("1011100100100110", '1', '1', "11", "010", "110", "001", '0', '-', "00"), -- i=1816
      ("1011100100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1817
      ("0101000100100000", '0', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1818
      ("0101100100100000", '1', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1819
      ("0101100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1820
      ("0100000100100000", '0', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1821
      ("0100100100100000", '1', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1822
      ("0100100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1823
      ("0000000110111001", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1824
      ("0000100110111001", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1825
      ("0000100110111001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1826
      ("1000000100100111", '0', '1', "00", "010", "111", "001", '0', '-', "00"), -- i=1827
      ("1000100100100111", '1', '1', "00", "010", "111", "001", '0', '-', "00"), -- i=1828
      ("1000100100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1829
      ("1001000100100111", '0', '1', "01", "010", "111", "001", '0', '-', "00"), -- i=1830
      ("1001100100100111", '1', '1', "01", "010", "111", "001", '0', '-', "00"), -- i=1831
      ("1001100100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1832
      ("1010000100100111", '0', '1', "10", "010", "111", "001", '0', '-', "00"), -- i=1833
      ("1010100100100111", '1', '1', "10", "010", "111", "001", '0', '-', "00"), -- i=1834
      ("1010100100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1835
      ("1011000100100111", '0', '1', "11", "010", "111", "001", '0', '-', "00"), -- i=1836
      ("1011100100100111", '1', '1', "11", "010", "111", "001", '0', '-', "00"), -- i=1837
      ("1011100100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1838
      ("0101000100100000", '0', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1839
      ("0101100100100000", '1', '1', "--", "010", "---", "001", '0', '1', "01"), -- i=1840
      ("0101100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1841
      ("0100000100100000", '0', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1842
      ("0100100100100000", '1', '0', "--", "010", "001", "---", '1', '-', "--"), -- i=1843
      ("0100100100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1844
      ("0000000111001100", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1845
      ("0000100111001100", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1846
      ("0000100111001100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1847
      ("1000000100110000", '0', '1', "00", "011", "000", "001", '0', '-', "00"), -- i=1848
      ("1000100100110000", '1', '1', "00", "011", "000", "001", '0', '-', "00"), -- i=1849
      ("1000100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1850
      ("1001000100110000", '0', '1', "01", "011", "000", "001", '0', '-', "00"), -- i=1851
      ("1001100100110000", '1', '1', "01", "011", "000", "001", '0', '-', "00"), -- i=1852
      ("1001100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1853
      ("1010000100110000", '0', '1', "10", "011", "000", "001", '0', '-', "00"), -- i=1854
      ("1010100100110000", '1', '1', "10", "011", "000", "001", '0', '-', "00"), -- i=1855
      ("1010100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1856
      ("1011000100110000", '0', '1', "11", "011", "000", "001", '0', '-', "00"), -- i=1857
      ("1011100100110000", '1', '1', "11", "011", "000", "001", '0', '-', "00"), -- i=1858
      ("1011100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1859
      ("0101000100110000", '0', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=1860
      ("0101100100110000", '1', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=1861
      ("0101100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1862
      ("0100000100110000", '0', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=1863
      ("0100100100110000", '1', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=1864
      ("0100100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1865
      ("0000000100100001", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1866
      ("0000100100100001", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1867
      ("0000100100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1868
      ("1000000100110001", '0', '1', "00", "011", "001", "001", '0', '-', "00"), -- i=1869
      ("1000100100110001", '1', '1', "00", "011", "001", "001", '0', '-', "00"), -- i=1870
      ("1000100100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1871
      ("1001000100110001", '0', '1', "01", "011", "001", "001", '0', '-', "00"), -- i=1872
      ("1001100100110001", '1', '1', "01", "011", "001", "001", '0', '-', "00"), -- i=1873
      ("1001100100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1874
      ("1010000100110001", '0', '1', "10", "011", "001", "001", '0', '-', "00"), -- i=1875
      ("1010100100110001", '1', '1', "10", "011", "001", "001", '0', '-', "00"), -- i=1876
      ("1010100100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1877
      ("1011000100110001", '0', '1', "11", "011", "001", "001", '0', '-', "00"), -- i=1878
      ("1011100100110001", '1', '1', "11", "011", "001", "001", '0', '-', "00"), -- i=1879
      ("1011100100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1880
      ("0101000100110000", '0', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=1881
      ("0101100100110000", '1', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=1882
      ("0101100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1883
      ("0100000100110000", '0', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=1884
      ("0100100100110000", '1', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=1885
      ("0100100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1886
      ("0000000111011010", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1887
      ("0000100111011010", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1888
      ("0000100111011010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1889
      ("1000000100110010", '0', '1', "00", "011", "010", "001", '0', '-', "00"), -- i=1890
      ("1000100100110010", '1', '1', "00", "011", "010", "001", '0', '-', "00"), -- i=1891
      ("1000100100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1892
      ("1001000100110010", '0', '1', "01", "011", "010", "001", '0', '-', "00"), -- i=1893
      ("1001100100110010", '1', '1', "01", "011", "010", "001", '0', '-', "00"), -- i=1894
      ("1001100100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1895
      ("1010000100110010", '0', '1', "10", "011", "010", "001", '0', '-', "00"), -- i=1896
      ("1010100100110010", '1', '1', "10", "011", "010", "001", '0', '-', "00"), -- i=1897
      ("1010100100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1898
      ("1011000100110010", '0', '1', "11", "011", "010", "001", '0', '-', "00"), -- i=1899
      ("1011100100110010", '1', '1', "11", "011", "010", "001", '0', '-', "00"), -- i=1900
      ("1011100100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1901
      ("0101000100110000", '0', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=1902
      ("0101100100110000", '1', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=1903
      ("0101100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1904
      ("0100000100110000", '0', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=1905
      ("0100100100110000", '1', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=1906
      ("0100100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1907
      ("0000000101010101", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1908
      ("0000100101010101", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1909
      ("0000100101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1910
      ("1000000100110011", '0', '1', "00", "011", "011", "001", '0', '-', "00"), -- i=1911
      ("1000100100110011", '1', '1', "00", "011", "011", "001", '0', '-', "00"), -- i=1912
      ("1000100100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1913
      ("1001000100110011", '0', '1', "01", "011", "011", "001", '0', '-', "00"), -- i=1914
      ("1001100100110011", '1', '1', "01", "011", "011", "001", '0', '-', "00"), -- i=1915
      ("1001100100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1916
      ("1010000100110011", '0', '1', "10", "011", "011", "001", '0', '-', "00"), -- i=1917
      ("1010100100110011", '1', '1', "10", "011", "011", "001", '0', '-', "00"), -- i=1918
      ("1010100100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1919
      ("1011000100110011", '0', '1', "11", "011", "011", "001", '0', '-', "00"), -- i=1920
      ("1011100100110011", '1', '1', "11", "011", "011", "001", '0', '-', "00"), -- i=1921
      ("1011100100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1922
      ("0101000100110000", '0', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=1923
      ("0101100100110000", '1', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=1924
      ("0101100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1925
      ("0100000100110000", '0', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=1926
      ("0100100100110000", '1', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=1927
      ("0100100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1928
      ("0000000111000011", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1929
      ("0000100111000011", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1930
      ("0000100111000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1931
      ("1000000100110100", '0', '1', "00", "011", "100", "001", '0', '-', "00"), -- i=1932
      ("1000100100110100", '1', '1', "00", "011", "100", "001", '0', '-', "00"), -- i=1933
      ("1000100100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1934
      ("1001000100110100", '0', '1', "01", "011", "100", "001", '0', '-', "00"), -- i=1935
      ("1001100100110100", '1', '1', "01", "011", "100", "001", '0', '-', "00"), -- i=1936
      ("1001100100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1937
      ("1010000100110100", '0', '1', "10", "011", "100", "001", '0', '-', "00"), -- i=1938
      ("1010100100110100", '1', '1', "10", "011", "100", "001", '0', '-', "00"), -- i=1939
      ("1010100100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1940
      ("1011000100110100", '0', '1', "11", "011", "100", "001", '0', '-', "00"), -- i=1941
      ("1011100100110100", '1', '1', "11", "011", "100", "001", '0', '-', "00"), -- i=1942
      ("1011100100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1943
      ("0101000100110000", '0', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=1944
      ("0101100100110000", '1', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=1945
      ("0101100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1946
      ("0100000100110000", '0', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=1947
      ("0100100100110000", '1', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=1948
      ("0100100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1949
      ("0000000101001011", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1950
      ("0000100101001011", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1951
      ("0000100101001011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1952
      ("1000000100110101", '0', '1', "00", "011", "101", "001", '0', '-', "00"), -- i=1953
      ("1000100100110101", '1', '1', "00", "011", "101", "001", '0', '-', "00"), -- i=1954
      ("1000100100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1955
      ("1001000100110101", '0', '1', "01", "011", "101", "001", '0', '-', "00"), -- i=1956
      ("1001100100110101", '1', '1', "01", "011", "101", "001", '0', '-', "00"), -- i=1957
      ("1001100100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1958
      ("1010000100110101", '0', '1', "10", "011", "101", "001", '0', '-', "00"), -- i=1959
      ("1010100100110101", '1', '1', "10", "011", "101", "001", '0', '-', "00"), -- i=1960
      ("1010100100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1961
      ("1011000100110101", '0', '1', "11", "011", "101", "001", '0', '-', "00"), -- i=1962
      ("1011100100110101", '1', '1', "11", "011", "101", "001", '0', '-', "00"), -- i=1963
      ("1011100100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1964
      ("0101000100110000", '0', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=1965
      ("0101100100110000", '1', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=1966
      ("0101100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1967
      ("0100000100110000", '0', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=1968
      ("0100100100110000", '1', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=1969
      ("0100100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1970
      ("0000000100011100", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1971
      ("0000100100011100", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1972
      ("0000100100011100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1973
      ("1000000100110110", '0', '1', "00", "011", "110", "001", '0', '-', "00"), -- i=1974
      ("1000100100110110", '1', '1', "00", "011", "110", "001", '0', '-', "00"), -- i=1975
      ("1000100100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1976
      ("1001000100110110", '0', '1', "01", "011", "110", "001", '0', '-', "00"), -- i=1977
      ("1001100100110110", '1', '1', "01", "011", "110", "001", '0', '-', "00"), -- i=1978
      ("1001100100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1979
      ("1010000100110110", '0', '1', "10", "011", "110", "001", '0', '-', "00"), -- i=1980
      ("1010100100110110", '1', '1', "10", "011", "110", "001", '0', '-', "00"), -- i=1981
      ("1010100100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1982
      ("1011000100110110", '0', '1', "11", "011", "110", "001", '0', '-', "00"), -- i=1983
      ("1011100100110110", '1', '1', "11", "011", "110", "001", '0', '-', "00"), -- i=1984
      ("1011100100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1985
      ("0101000100110000", '0', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=1986
      ("0101100100110000", '1', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=1987
      ("0101100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1988
      ("0100000100110000", '0', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=1989
      ("0100100100110000", '1', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=1990
      ("0100100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1991
      ("0000000101011100", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1992
      ("0000100101011100", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=1993
      ("0000100101011100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1994
      ("1000000100110111", '0', '1', "00", "011", "111", "001", '0', '-', "00"), -- i=1995
      ("1000100100110111", '1', '1', "00", "011", "111", "001", '0', '-', "00"), -- i=1996
      ("1000100100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=1997
      ("1001000100110111", '0', '1', "01", "011", "111", "001", '0', '-', "00"), -- i=1998
      ("1001100100110111", '1', '1', "01", "011", "111", "001", '0', '-', "00"), -- i=1999
      ("1001100100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2000
      ("1010000100110111", '0', '1', "10", "011", "111", "001", '0', '-', "00"), -- i=2001
      ("1010100100110111", '1', '1', "10", "011", "111", "001", '0', '-', "00"), -- i=2002
      ("1010100100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2003
      ("1011000100110111", '0', '1', "11", "011", "111", "001", '0', '-', "00"), -- i=2004
      ("1011100100110111", '1', '1', "11", "011", "111", "001", '0', '-', "00"), -- i=2005
      ("1011100100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2006
      ("0101000100110000", '0', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=2007
      ("0101100100110000", '1', '1', "--", "011", "---", "001", '0', '1', "01"), -- i=2008
      ("0101100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2009
      ("0100000100110000", '0', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=2010
      ("0100100100110000", '1', '0', "--", "011", "001", "---", '1', '-', "--"), -- i=2011
      ("0100100100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2012
      ("0000000111000110", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2013
      ("0000100111000110", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2014
      ("0000100111000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2015
      ("1000000101000000", '0', '1', "00", "100", "000", "001", '0', '-', "00"), -- i=2016
      ("1000100101000000", '1', '1', "00", "100", "000", "001", '0', '-', "00"), -- i=2017
      ("1000100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2018
      ("1001000101000000", '0', '1', "01", "100", "000", "001", '0', '-', "00"), -- i=2019
      ("1001100101000000", '1', '1', "01", "100", "000", "001", '0', '-', "00"), -- i=2020
      ("1001100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2021
      ("1010000101000000", '0', '1', "10", "100", "000", "001", '0', '-', "00"), -- i=2022
      ("1010100101000000", '1', '1', "10", "100", "000", "001", '0', '-', "00"), -- i=2023
      ("1010100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2024
      ("1011000101000000", '0', '1', "11", "100", "000", "001", '0', '-', "00"), -- i=2025
      ("1011100101000000", '1', '1', "11", "100", "000", "001", '0', '-', "00"), -- i=2026
      ("1011100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2027
      ("0101000101000000", '0', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2028
      ("0101100101000000", '1', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2029
      ("0101100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2030
      ("0100000101000000", '0', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2031
      ("0100100101000000", '1', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2032
      ("0100100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2033
      ("0000000100000100", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2034
      ("0000100100000100", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2035
      ("0000100100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2036
      ("1000000101000001", '0', '1', "00", "100", "001", "001", '0', '-', "00"), -- i=2037
      ("1000100101000001", '1', '1', "00", "100", "001", "001", '0', '-', "00"), -- i=2038
      ("1000100101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2039
      ("1001000101000001", '0', '1', "01", "100", "001", "001", '0', '-', "00"), -- i=2040
      ("1001100101000001", '1', '1', "01", "100", "001", "001", '0', '-', "00"), -- i=2041
      ("1001100101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2042
      ("1010000101000001", '0', '1', "10", "100", "001", "001", '0', '-', "00"), -- i=2043
      ("1010100101000001", '1', '1', "10", "100", "001", "001", '0', '-', "00"), -- i=2044
      ("1010100101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2045
      ("1011000101000001", '0', '1', "11", "100", "001", "001", '0', '-', "00"), -- i=2046
      ("1011100101000001", '1', '1', "11", "100", "001", "001", '0', '-', "00"), -- i=2047
      ("1011100101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2048
      ("0101000101000000", '0', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2049
      ("0101100101000000", '1', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2050
      ("0101100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2051
      ("0100000101000000", '0', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2052
      ("0100100101000000", '1', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2053
      ("0100100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2054
      ("0000000110000011", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2055
      ("0000100110000011", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2056
      ("0000100110000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2057
      ("1000000101000010", '0', '1', "00", "100", "010", "001", '0', '-', "00"), -- i=2058
      ("1000100101000010", '1', '1', "00", "100", "010", "001", '0', '-', "00"), -- i=2059
      ("1000100101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2060
      ("1001000101000010", '0', '1', "01", "100", "010", "001", '0', '-', "00"), -- i=2061
      ("1001100101000010", '1', '1', "01", "100", "010", "001", '0', '-', "00"), -- i=2062
      ("1001100101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2063
      ("1010000101000010", '0', '1', "10", "100", "010", "001", '0', '-', "00"), -- i=2064
      ("1010100101000010", '1', '1', "10", "100", "010", "001", '0', '-', "00"), -- i=2065
      ("1010100101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2066
      ("1011000101000010", '0', '1', "11", "100", "010", "001", '0', '-', "00"), -- i=2067
      ("1011100101000010", '1', '1', "11", "100", "010", "001", '0', '-', "00"), -- i=2068
      ("1011100101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2069
      ("0101000101000000", '0', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2070
      ("0101100101000000", '1', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2071
      ("0101100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2072
      ("0100000101000000", '0', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2073
      ("0100100101000000", '1', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2074
      ("0100100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2075
      ("0000000110011011", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2076
      ("0000100110011011", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2077
      ("0000100110011011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2078
      ("1000000101000011", '0', '1', "00", "100", "011", "001", '0', '-', "00"), -- i=2079
      ("1000100101000011", '1', '1', "00", "100", "011", "001", '0', '-', "00"), -- i=2080
      ("1000100101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2081
      ("1001000101000011", '0', '1', "01", "100", "011", "001", '0', '-', "00"), -- i=2082
      ("1001100101000011", '1', '1', "01", "100", "011", "001", '0', '-', "00"), -- i=2083
      ("1001100101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2084
      ("1010000101000011", '0', '1', "10", "100", "011", "001", '0', '-', "00"), -- i=2085
      ("1010100101000011", '1', '1', "10", "100", "011", "001", '0', '-', "00"), -- i=2086
      ("1010100101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2087
      ("1011000101000011", '0', '1', "11", "100", "011", "001", '0', '-', "00"), -- i=2088
      ("1011100101000011", '1', '1', "11", "100", "011", "001", '0', '-', "00"), -- i=2089
      ("1011100101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2090
      ("0101000101000000", '0', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2091
      ("0101100101000000", '1', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2092
      ("0101100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2093
      ("0100000101000000", '0', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2094
      ("0100100101000000", '1', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2095
      ("0100100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2096
      ("0000000101000111", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2097
      ("0000100101000111", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2098
      ("0000100101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2099
      ("1000000101000100", '0', '1', "00", "100", "100", "001", '0', '-', "00"), -- i=2100
      ("1000100101000100", '1', '1', "00", "100", "100", "001", '0', '-', "00"), -- i=2101
      ("1000100101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2102
      ("1001000101000100", '0', '1', "01", "100", "100", "001", '0', '-', "00"), -- i=2103
      ("1001100101000100", '1', '1', "01", "100", "100", "001", '0', '-', "00"), -- i=2104
      ("1001100101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2105
      ("1010000101000100", '0', '1', "10", "100", "100", "001", '0', '-', "00"), -- i=2106
      ("1010100101000100", '1', '1', "10", "100", "100", "001", '0', '-', "00"), -- i=2107
      ("1010100101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2108
      ("1011000101000100", '0', '1', "11", "100", "100", "001", '0', '-', "00"), -- i=2109
      ("1011100101000100", '1', '1', "11", "100", "100", "001", '0', '-', "00"), -- i=2110
      ("1011100101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2111
      ("0101000101000000", '0', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2112
      ("0101100101000000", '1', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2113
      ("0101100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2114
      ("0100000101000000", '0', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2115
      ("0100100101000000", '1', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2116
      ("0100100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2117
      ("0000000111011011", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2118
      ("0000100111011011", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2119
      ("0000100111011011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2120
      ("1000000101000101", '0', '1', "00", "100", "101", "001", '0', '-', "00"), -- i=2121
      ("1000100101000101", '1', '1', "00", "100", "101", "001", '0', '-', "00"), -- i=2122
      ("1000100101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2123
      ("1001000101000101", '0', '1', "01", "100", "101", "001", '0', '-', "00"), -- i=2124
      ("1001100101000101", '1', '1', "01", "100", "101", "001", '0', '-', "00"), -- i=2125
      ("1001100101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2126
      ("1010000101000101", '0', '1', "10", "100", "101", "001", '0', '-', "00"), -- i=2127
      ("1010100101000101", '1', '1', "10", "100", "101", "001", '0', '-', "00"), -- i=2128
      ("1010100101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2129
      ("1011000101000101", '0', '1', "11", "100", "101", "001", '0', '-', "00"), -- i=2130
      ("1011100101000101", '1', '1', "11", "100", "101", "001", '0', '-', "00"), -- i=2131
      ("1011100101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2132
      ("0101000101000000", '0', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2133
      ("0101100101000000", '1', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2134
      ("0101100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2135
      ("0100000101000000", '0', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2136
      ("0100100101000000", '1', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2137
      ("0100100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2138
      ("0000000100001000", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2139
      ("0000100100001000", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2140
      ("0000100100001000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2141
      ("1000000101000110", '0', '1', "00", "100", "110", "001", '0', '-', "00"), -- i=2142
      ("1000100101000110", '1', '1', "00", "100", "110", "001", '0', '-', "00"), -- i=2143
      ("1000100101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2144
      ("1001000101000110", '0', '1', "01", "100", "110", "001", '0', '-', "00"), -- i=2145
      ("1001100101000110", '1', '1', "01", "100", "110", "001", '0', '-', "00"), -- i=2146
      ("1001100101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2147
      ("1010000101000110", '0', '1', "10", "100", "110", "001", '0', '-', "00"), -- i=2148
      ("1010100101000110", '1', '1', "10", "100", "110", "001", '0', '-', "00"), -- i=2149
      ("1010100101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2150
      ("1011000101000110", '0', '1', "11", "100", "110", "001", '0', '-', "00"), -- i=2151
      ("1011100101000110", '1', '1', "11", "100", "110", "001", '0', '-', "00"), -- i=2152
      ("1011100101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2153
      ("0101000101000000", '0', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2154
      ("0101100101000000", '1', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2155
      ("0101100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2156
      ("0100000101000000", '0', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2157
      ("0100100101000000", '1', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2158
      ("0100100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2159
      ("0000000111011111", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2160
      ("0000100111011111", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2161
      ("0000100111011111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2162
      ("1000000101000111", '0', '1', "00", "100", "111", "001", '0', '-', "00"), -- i=2163
      ("1000100101000111", '1', '1', "00", "100", "111", "001", '0', '-', "00"), -- i=2164
      ("1000100101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2165
      ("1001000101000111", '0', '1', "01", "100", "111", "001", '0', '-', "00"), -- i=2166
      ("1001100101000111", '1', '1', "01", "100", "111", "001", '0', '-', "00"), -- i=2167
      ("1001100101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2168
      ("1010000101000111", '0', '1', "10", "100", "111", "001", '0', '-', "00"), -- i=2169
      ("1010100101000111", '1', '1', "10", "100", "111", "001", '0', '-', "00"), -- i=2170
      ("1010100101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2171
      ("1011000101000111", '0', '1', "11", "100", "111", "001", '0', '-', "00"), -- i=2172
      ("1011100101000111", '1', '1', "11", "100", "111", "001", '0', '-', "00"), -- i=2173
      ("1011100101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2174
      ("0101000101000000", '0', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2175
      ("0101100101000000", '1', '1', "--", "100", "---", "001", '0', '1', "01"), -- i=2176
      ("0101100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2177
      ("0100000101000000", '0', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2178
      ("0100100101000000", '1', '0', "--", "100", "001", "---", '1', '-', "--"), -- i=2179
      ("0100100101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2180
      ("0000000100100100", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2181
      ("0000100100100100", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2182
      ("0000100100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2183
      ("1000000101010000", '0', '1', "00", "101", "000", "001", '0', '-', "00"), -- i=2184
      ("1000100101010000", '1', '1', "00", "101", "000", "001", '0', '-', "00"), -- i=2185
      ("1000100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2186
      ("1001000101010000", '0', '1', "01", "101", "000", "001", '0', '-', "00"), -- i=2187
      ("1001100101010000", '1', '1', "01", "101", "000", "001", '0', '-', "00"), -- i=2188
      ("1001100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2189
      ("1010000101010000", '0', '1', "10", "101", "000", "001", '0', '-', "00"), -- i=2190
      ("1010100101010000", '1', '1', "10", "101", "000", "001", '0', '-', "00"), -- i=2191
      ("1010100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2192
      ("1011000101010000", '0', '1', "11", "101", "000", "001", '0', '-', "00"), -- i=2193
      ("1011100101010000", '1', '1', "11", "101", "000", "001", '0', '-', "00"), -- i=2194
      ("1011100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2195
      ("0101000101010000", '0', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2196
      ("0101100101010000", '1', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2197
      ("0101100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2198
      ("0100000101010000", '0', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2199
      ("0100100101010000", '1', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2200
      ("0100100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2201
      ("0000000100001100", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2202
      ("0000100100001100", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2203
      ("0000100100001100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2204
      ("1000000101010001", '0', '1', "00", "101", "001", "001", '0', '-', "00"), -- i=2205
      ("1000100101010001", '1', '1', "00", "101", "001", "001", '0', '-', "00"), -- i=2206
      ("1000100101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2207
      ("1001000101010001", '0', '1', "01", "101", "001", "001", '0', '-', "00"), -- i=2208
      ("1001100101010001", '1', '1', "01", "101", "001", "001", '0', '-', "00"), -- i=2209
      ("1001100101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2210
      ("1010000101010001", '0', '1', "10", "101", "001", "001", '0', '-', "00"), -- i=2211
      ("1010100101010001", '1', '1', "10", "101", "001", "001", '0', '-', "00"), -- i=2212
      ("1010100101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2213
      ("1011000101010001", '0', '1', "11", "101", "001", "001", '0', '-', "00"), -- i=2214
      ("1011100101010001", '1', '1', "11", "101", "001", "001", '0', '-', "00"), -- i=2215
      ("1011100101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2216
      ("0101000101010000", '0', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2217
      ("0101100101010000", '1', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2218
      ("0101100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2219
      ("0100000101010000", '0', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2220
      ("0100100101010000", '1', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2221
      ("0100100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2222
      ("0000000110000000", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2223
      ("0000100110000000", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2224
      ("0000100110000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2225
      ("1000000101010010", '0', '1', "00", "101", "010", "001", '0', '-', "00"), -- i=2226
      ("1000100101010010", '1', '1', "00", "101", "010", "001", '0', '-', "00"), -- i=2227
      ("1000100101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2228
      ("1001000101010010", '0', '1', "01", "101", "010", "001", '0', '-', "00"), -- i=2229
      ("1001100101010010", '1', '1', "01", "101", "010", "001", '0', '-', "00"), -- i=2230
      ("1001100101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2231
      ("1010000101010010", '0', '1', "10", "101", "010", "001", '0', '-', "00"), -- i=2232
      ("1010100101010010", '1', '1', "10", "101", "010", "001", '0', '-', "00"), -- i=2233
      ("1010100101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2234
      ("1011000101010010", '0', '1', "11", "101", "010", "001", '0', '-', "00"), -- i=2235
      ("1011100101010010", '1', '1', "11", "101", "010", "001", '0', '-', "00"), -- i=2236
      ("1011100101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2237
      ("0101000101010000", '0', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2238
      ("0101100101010000", '1', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2239
      ("0101100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2240
      ("0100000101010000", '0', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2241
      ("0100100101010000", '1', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2242
      ("0100100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2243
      ("0000000111110011", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2244
      ("0000100111110011", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2245
      ("0000100111110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2246
      ("1000000101010011", '0', '1', "00", "101", "011", "001", '0', '-', "00"), -- i=2247
      ("1000100101010011", '1', '1', "00", "101", "011", "001", '0', '-', "00"), -- i=2248
      ("1000100101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2249
      ("1001000101010011", '0', '1', "01", "101", "011", "001", '0', '-', "00"), -- i=2250
      ("1001100101010011", '1', '1', "01", "101", "011", "001", '0', '-', "00"), -- i=2251
      ("1001100101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2252
      ("1010000101010011", '0', '1', "10", "101", "011", "001", '0', '-', "00"), -- i=2253
      ("1010100101010011", '1', '1', "10", "101", "011", "001", '0', '-', "00"), -- i=2254
      ("1010100101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2255
      ("1011000101010011", '0', '1', "11", "101", "011", "001", '0', '-', "00"), -- i=2256
      ("1011100101010011", '1', '1', "11", "101", "011", "001", '0', '-', "00"), -- i=2257
      ("1011100101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2258
      ("0101000101010000", '0', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2259
      ("0101100101010000", '1', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2260
      ("0101100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2261
      ("0100000101010000", '0', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2262
      ("0100100101010000", '1', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2263
      ("0100100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2264
      ("0000000111011001", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2265
      ("0000100111011001", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2266
      ("0000100111011001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2267
      ("1000000101010100", '0', '1', "00", "101", "100", "001", '0', '-', "00"), -- i=2268
      ("1000100101010100", '1', '1', "00", "101", "100", "001", '0', '-', "00"), -- i=2269
      ("1000100101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2270
      ("1001000101010100", '0', '1', "01", "101", "100", "001", '0', '-', "00"), -- i=2271
      ("1001100101010100", '1', '1', "01", "101", "100", "001", '0', '-', "00"), -- i=2272
      ("1001100101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2273
      ("1010000101010100", '0', '1', "10", "101", "100", "001", '0', '-', "00"), -- i=2274
      ("1010100101010100", '1', '1', "10", "101", "100", "001", '0', '-', "00"), -- i=2275
      ("1010100101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2276
      ("1011000101010100", '0', '1', "11", "101", "100", "001", '0', '-', "00"), -- i=2277
      ("1011100101010100", '1', '1', "11", "101", "100", "001", '0', '-', "00"), -- i=2278
      ("1011100101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2279
      ("0101000101010000", '0', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2280
      ("0101100101010000", '1', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2281
      ("0101100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2282
      ("0100000101010000", '0', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2283
      ("0100100101010000", '1', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2284
      ("0100100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2285
      ("0000000100110101", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2286
      ("0000100100110101", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2287
      ("0000100100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2288
      ("1000000101010101", '0', '1', "00", "101", "101", "001", '0', '-', "00"), -- i=2289
      ("1000100101010101", '1', '1', "00", "101", "101", "001", '0', '-', "00"), -- i=2290
      ("1000100101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2291
      ("1001000101010101", '0', '1', "01", "101", "101", "001", '0', '-', "00"), -- i=2292
      ("1001100101010101", '1', '1', "01", "101", "101", "001", '0', '-', "00"), -- i=2293
      ("1001100101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2294
      ("1010000101010101", '0', '1', "10", "101", "101", "001", '0', '-', "00"), -- i=2295
      ("1010100101010101", '1', '1', "10", "101", "101", "001", '0', '-', "00"), -- i=2296
      ("1010100101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2297
      ("1011000101010101", '0', '1', "11", "101", "101", "001", '0', '-', "00"), -- i=2298
      ("1011100101010101", '1', '1', "11", "101", "101", "001", '0', '-', "00"), -- i=2299
      ("1011100101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2300
      ("0101000101010000", '0', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2301
      ("0101100101010000", '1', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2302
      ("0101100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2303
      ("0100000101010000", '0', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2304
      ("0100100101010000", '1', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2305
      ("0100100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2306
      ("0000000100100111", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2307
      ("0000100100100111", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2308
      ("0000100100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2309
      ("1000000101010110", '0', '1', "00", "101", "110", "001", '0', '-', "00"), -- i=2310
      ("1000100101010110", '1', '1', "00", "101", "110", "001", '0', '-', "00"), -- i=2311
      ("1000100101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2312
      ("1001000101010110", '0', '1', "01", "101", "110", "001", '0', '-', "00"), -- i=2313
      ("1001100101010110", '1', '1', "01", "101", "110", "001", '0', '-', "00"), -- i=2314
      ("1001100101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2315
      ("1010000101010110", '0', '1', "10", "101", "110", "001", '0', '-', "00"), -- i=2316
      ("1010100101010110", '1', '1', "10", "101", "110", "001", '0', '-', "00"), -- i=2317
      ("1010100101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2318
      ("1011000101010110", '0', '1', "11", "101", "110", "001", '0', '-', "00"), -- i=2319
      ("1011100101010110", '1', '1', "11", "101", "110", "001", '0', '-', "00"), -- i=2320
      ("1011100101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2321
      ("0101000101010000", '0', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2322
      ("0101100101010000", '1', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2323
      ("0101100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2324
      ("0100000101010000", '0', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2325
      ("0100100101010000", '1', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2326
      ("0100100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2327
      ("0000000101010010", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2328
      ("0000100101010010", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2329
      ("0000100101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2330
      ("1000000101010111", '0', '1', "00", "101", "111", "001", '0', '-', "00"), -- i=2331
      ("1000100101010111", '1', '1', "00", "101", "111", "001", '0', '-', "00"), -- i=2332
      ("1000100101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2333
      ("1001000101010111", '0', '1', "01", "101", "111", "001", '0', '-', "00"), -- i=2334
      ("1001100101010111", '1', '1', "01", "101", "111", "001", '0', '-', "00"), -- i=2335
      ("1001100101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2336
      ("1010000101010111", '0', '1', "10", "101", "111", "001", '0', '-', "00"), -- i=2337
      ("1010100101010111", '1', '1', "10", "101", "111", "001", '0', '-', "00"), -- i=2338
      ("1010100101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2339
      ("1011000101010111", '0', '1', "11", "101", "111", "001", '0', '-', "00"), -- i=2340
      ("1011100101010111", '1', '1', "11", "101", "111", "001", '0', '-', "00"), -- i=2341
      ("1011100101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2342
      ("0101000101010000", '0', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2343
      ("0101100101010000", '1', '1', "--", "101", "---", "001", '0', '1', "01"), -- i=2344
      ("0101100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2345
      ("0100000101010000", '0', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2346
      ("0100100101010000", '1', '0', "--", "101", "001", "---", '1', '-', "--"), -- i=2347
      ("0100100101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2348
      ("0000000110001010", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2349
      ("0000100110001010", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2350
      ("0000100110001010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2351
      ("1000000101100000", '0', '1', "00", "110", "000", "001", '0', '-', "00"), -- i=2352
      ("1000100101100000", '1', '1', "00", "110", "000", "001", '0', '-', "00"), -- i=2353
      ("1000100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2354
      ("1001000101100000", '0', '1', "01", "110", "000", "001", '0', '-', "00"), -- i=2355
      ("1001100101100000", '1', '1', "01", "110", "000", "001", '0', '-', "00"), -- i=2356
      ("1001100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2357
      ("1010000101100000", '0', '1', "10", "110", "000", "001", '0', '-', "00"), -- i=2358
      ("1010100101100000", '1', '1', "10", "110", "000", "001", '0', '-', "00"), -- i=2359
      ("1010100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2360
      ("1011000101100000", '0', '1', "11", "110", "000", "001", '0', '-', "00"), -- i=2361
      ("1011100101100000", '1', '1', "11", "110", "000", "001", '0', '-', "00"), -- i=2362
      ("1011100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2363
      ("0101000101100000", '0', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2364
      ("0101100101100000", '1', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2365
      ("0101100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2366
      ("0100000101100000", '0', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2367
      ("0100100101100000", '1', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2368
      ("0100100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2369
      ("0000000111010101", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2370
      ("0000100111010101", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2371
      ("0000100111010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2372
      ("1000000101100001", '0', '1', "00", "110", "001", "001", '0', '-', "00"), -- i=2373
      ("1000100101100001", '1', '1', "00", "110", "001", "001", '0', '-', "00"), -- i=2374
      ("1000100101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2375
      ("1001000101100001", '0', '1', "01", "110", "001", "001", '0', '-', "00"), -- i=2376
      ("1001100101100001", '1', '1', "01", "110", "001", "001", '0', '-', "00"), -- i=2377
      ("1001100101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2378
      ("1010000101100001", '0', '1', "10", "110", "001", "001", '0', '-', "00"), -- i=2379
      ("1010100101100001", '1', '1', "10", "110", "001", "001", '0', '-', "00"), -- i=2380
      ("1010100101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2381
      ("1011000101100001", '0', '1', "11", "110", "001", "001", '0', '-', "00"), -- i=2382
      ("1011100101100001", '1', '1', "11", "110", "001", "001", '0', '-', "00"), -- i=2383
      ("1011100101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2384
      ("0101000101100000", '0', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2385
      ("0101100101100000", '1', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2386
      ("0101100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2387
      ("0100000101100000", '0', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2388
      ("0100100101100000", '1', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2389
      ("0100100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2390
      ("0000000100011011", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2391
      ("0000100100011011", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2392
      ("0000100100011011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2393
      ("1000000101100010", '0', '1', "00", "110", "010", "001", '0', '-', "00"), -- i=2394
      ("1000100101100010", '1', '1', "00", "110", "010", "001", '0', '-', "00"), -- i=2395
      ("1000100101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2396
      ("1001000101100010", '0', '1', "01", "110", "010", "001", '0', '-', "00"), -- i=2397
      ("1001100101100010", '1', '1', "01", "110", "010", "001", '0', '-', "00"), -- i=2398
      ("1001100101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2399
      ("1010000101100010", '0', '1', "10", "110", "010", "001", '0', '-', "00"), -- i=2400
      ("1010100101100010", '1', '1', "10", "110", "010", "001", '0', '-', "00"), -- i=2401
      ("1010100101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2402
      ("1011000101100010", '0', '1', "11", "110", "010", "001", '0', '-', "00"), -- i=2403
      ("1011100101100010", '1', '1', "11", "110", "010", "001", '0', '-', "00"), -- i=2404
      ("1011100101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2405
      ("0101000101100000", '0', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2406
      ("0101100101100000", '1', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2407
      ("0101100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2408
      ("0100000101100000", '0', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2409
      ("0100100101100000", '1', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2410
      ("0100100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2411
      ("0000000100011010", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2412
      ("0000100100011010", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2413
      ("0000100100011010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2414
      ("1000000101100011", '0', '1', "00", "110", "011", "001", '0', '-', "00"), -- i=2415
      ("1000100101100011", '1', '1', "00", "110", "011", "001", '0', '-', "00"), -- i=2416
      ("1000100101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2417
      ("1001000101100011", '0', '1', "01", "110", "011", "001", '0', '-', "00"), -- i=2418
      ("1001100101100011", '1', '1', "01", "110", "011", "001", '0', '-', "00"), -- i=2419
      ("1001100101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2420
      ("1010000101100011", '0', '1', "10", "110", "011", "001", '0', '-', "00"), -- i=2421
      ("1010100101100011", '1', '1', "10", "110", "011", "001", '0', '-', "00"), -- i=2422
      ("1010100101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2423
      ("1011000101100011", '0', '1', "11", "110", "011", "001", '0', '-', "00"), -- i=2424
      ("1011100101100011", '1', '1', "11", "110", "011", "001", '0', '-', "00"), -- i=2425
      ("1011100101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2426
      ("0101000101100000", '0', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2427
      ("0101100101100000", '1', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2428
      ("0101100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2429
      ("0100000101100000", '0', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2430
      ("0100100101100000", '1', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2431
      ("0100100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2432
      ("0000000100100101", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2433
      ("0000100100100101", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2434
      ("0000100100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2435
      ("1000000101100100", '0', '1', "00", "110", "100", "001", '0', '-', "00"), -- i=2436
      ("1000100101100100", '1', '1', "00", "110", "100", "001", '0', '-', "00"), -- i=2437
      ("1000100101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2438
      ("1001000101100100", '0', '1', "01", "110", "100", "001", '0', '-', "00"), -- i=2439
      ("1001100101100100", '1', '1', "01", "110", "100", "001", '0', '-', "00"), -- i=2440
      ("1001100101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2441
      ("1010000101100100", '0', '1', "10", "110", "100", "001", '0', '-', "00"), -- i=2442
      ("1010100101100100", '1', '1', "10", "110", "100", "001", '0', '-', "00"), -- i=2443
      ("1010100101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2444
      ("1011000101100100", '0', '1', "11", "110", "100", "001", '0', '-', "00"), -- i=2445
      ("1011100101100100", '1', '1', "11", "110", "100", "001", '0', '-', "00"), -- i=2446
      ("1011100101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2447
      ("0101000101100000", '0', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2448
      ("0101100101100000", '1', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2449
      ("0101100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2450
      ("0100000101100000", '0', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2451
      ("0100100101100000", '1', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2452
      ("0100100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2453
      ("0000000111000101", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2454
      ("0000100111000101", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2455
      ("0000100111000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2456
      ("1000000101100101", '0', '1', "00", "110", "101", "001", '0', '-', "00"), -- i=2457
      ("1000100101100101", '1', '1', "00", "110", "101", "001", '0', '-', "00"), -- i=2458
      ("1000100101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2459
      ("1001000101100101", '0', '1', "01", "110", "101", "001", '0', '-', "00"), -- i=2460
      ("1001100101100101", '1', '1', "01", "110", "101", "001", '0', '-', "00"), -- i=2461
      ("1001100101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2462
      ("1010000101100101", '0', '1', "10", "110", "101", "001", '0', '-', "00"), -- i=2463
      ("1010100101100101", '1', '1', "10", "110", "101", "001", '0', '-', "00"), -- i=2464
      ("1010100101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2465
      ("1011000101100101", '0', '1', "11", "110", "101", "001", '0', '-', "00"), -- i=2466
      ("1011100101100101", '1', '1', "11", "110", "101", "001", '0', '-', "00"), -- i=2467
      ("1011100101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2468
      ("0101000101100000", '0', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2469
      ("0101100101100000", '1', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2470
      ("0101100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2471
      ("0100000101100000", '0', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2472
      ("0100100101100000", '1', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2473
      ("0100100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2474
      ("0000000110111011", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2475
      ("0000100110111011", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2476
      ("0000100110111011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2477
      ("1000000101100110", '0', '1', "00", "110", "110", "001", '0', '-', "00"), -- i=2478
      ("1000100101100110", '1', '1', "00", "110", "110", "001", '0', '-', "00"), -- i=2479
      ("1000100101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2480
      ("1001000101100110", '0', '1', "01", "110", "110", "001", '0', '-', "00"), -- i=2481
      ("1001100101100110", '1', '1', "01", "110", "110", "001", '0', '-', "00"), -- i=2482
      ("1001100101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2483
      ("1010000101100110", '0', '1', "10", "110", "110", "001", '0', '-', "00"), -- i=2484
      ("1010100101100110", '1', '1', "10", "110", "110", "001", '0', '-', "00"), -- i=2485
      ("1010100101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2486
      ("1011000101100110", '0', '1', "11", "110", "110", "001", '0', '-', "00"), -- i=2487
      ("1011100101100110", '1', '1', "11", "110", "110", "001", '0', '-', "00"), -- i=2488
      ("1011100101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2489
      ("0101000101100000", '0', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2490
      ("0101100101100000", '1', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2491
      ("0101100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2492
      ("0100000101100000", '0', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2493
      ("0100100101100000", '1', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2494
      ("0100100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2495
      ("0000000100101110", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2496
      ("0000100100101110", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2497
      ("0000100100101110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2498
      ("1000000101100111", '0', '1', "00", "110", "111", "001", '0', '-', "00"), -- i=2499
      ("1000100101100111", '1', '1', "00", "110", "111", "001", '0', '-', "00"), -- i=2500
      ("1000100101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2501
      ("1001000101100111", '0', '1', "01", "110", "111", "001", '0', '-', "00"), -- i=2502
      ("1001100101100111", '1', '1', "01", "110", "111", "001", '0', '-', "00"), -- i=2503
      ("1001100101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2504
      ("1010000101100111", '0', '1', "10", "110", "111", "001", '0', '-', "00"), -- i=2505
      ("1010100101100111", '1', '1', "10", "110", "111", "001", '0', '-', "00"), -- i=2506
      ("1010100101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2507
      ("1011000101100111", '0', '1', "11", "110", "111", "001", '0', '-', "00"), -- i=2508
      ("1011100101100111", '1', '1', "11", "110", "111", "001", '0', '-', "00"), -- i=2509
      ("1011100101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2510
      ("0101000101100000", '0', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2511
      ("0101100101100000", '1', '1', "--", "110", "---", "001", '0', '1', "01"), -- i=2512
      ("0101100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2513
      ("0100000101100000", '0', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2514
      ("0100100101100000", '1', '0', "--", "110", "001", "---", '1', '-', "--"), -- i=2515
      ("0100100101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2516
      ("0000000100000000", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2517
      ("0000100100000000", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2518
      ("0000100100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2519
      ("1000000101110000", '0', '1', "00", "111", "000", "001", '0', '-', "00"), -- i=2520
      ("1000100101110000", '1', '1', "00", "111", "000", "001", '0', '-', "00"), -- i=2521
      ("1000100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2522
      ("1001000101110000", '0', '1', "01", "111", "000", "001", '0', '-', "00"), -- i=2523
      ("1001100101110000", '1', '1', "01", "111", "000", "001", '0', '-', "00"), -- i=2524
      ("1001100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2525
      ("1010000101110000", '0', '1', "10", "111", "000", "001", '0', '-', "00"), -- i=2526
      ("1010100101110000", '1', '1', "10", "111", "000", "001", '0', '-', "00"), -- i=2527
      ("1010100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2528
      ("1011000101110000", '0', '1', "11", "111", "000", "001", '0', '-', "00"), -- i=2529
      ("1011100101110000", '1', '1', "11", "111", "000", "001", '0', '-', "00"), -- i=2530
      ("1011100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2531
      ("0101000101110000", '0', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2532
      ("0101100101110000", '1', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2533
      ("0101100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2534
      ("0100000101110000", '0', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2535
      ("0100100101110000", '1', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2536
      ("0100100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2537
      ("0000000100000110", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2538
      ("0000100100000110", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2539
      ("0000100100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2540
      ("1000000101110001", '0', '1', "00", "111", "001", "001", '0', '-', "00"), -- i=2541
      ("1000100101110001", '1', '1', "00", "111", "001", "001", '0', '-', "00"), -- i=2542
      ("1000100101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2543
      ("1001000101110001", '0', '1', "01", "111", "001", "001", '0', '-', "00"), -- i=2544
      ("1001100101110001", '1', '1', "01", "111", "001", "001", '0', '-', "00"), -- i=2545
      ("1001100101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2546
      ("1010000101110001", '0', '1', "10", "111", "001", "001", '0', '-', "00"), -- i=2547
      ("1010100101110001", '1', '1', "10", "111", "001", "001", '0', '-', "00"), -- i=2548
      ("1010100101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2549
      ("1011000101110001", '0', '1', "11", "111", "001", "001", '0', '-', "00"), -- i=2550
      ("1011100101110001", '1', '1', "11", "111", "001", "001", '0', '-', "00"), -- i=2551
      ("1011100101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2552
      ("0101000101110000", '0', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2553
      ("0101100101110000", '1', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2554
      ("0101100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2555
      ("0100000101110000", '0', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2556
      ("0100100101110000", '1', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2557
      ("0100100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2558
      ("0000000110000110", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2559
      ("0000100110000110", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2560
      ("0000100110000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2561
      ("1000000101110010", '0', '1', "00", "111", "010", "001", '0', '-', "00"), -- i=2562
      ("1000100101110010", '1', '1', "00", "111", "010", "001", '0', '-', "00"), -- i=2563
      ("1000100101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2564
      ("1001000101110010", '0', '1', "01", "111", "010", "001", '0', '-', "00"), -- i=2565
      ("1001100101110010", '1', '1', "01", "111", "010", "001", '0', '-', "00"), -- i=2566
      ("1001100101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2567
      ("1010000101110010", '0', '1', "10", "111", "010", "001", '0', '-', "00"), -- i=2568
      ("1010100101110010", '1', '1', "10", "111", "010", "001", '0', '-', "00"), -- i=2569
      ("1010100101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2570
      ("1011000101110010", '0', '1', "11", "111", "010", "001", '0', '-', "00"), -- i=2571
      ("1011100101110010", '1', '1', "11", "111", "010", "001", '0', '-', "00"), -- i=2572
      ("1011100101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2573
      ("0101000101110000", '0', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2574
      ("0101100101110000", '1', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2575
      ("0101100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2576
      ("0100000101110000", '0', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2577
      ("0100100101110000", '1', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2578
      ("0100100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2579
      ("0000000111111110", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2580
      ("0000100111111110", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2581
      ("0000100111111110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2582
      ("1000000101110011", '0', '1', "00", "111", "011", "001", '0', '-', "00"), -- i=2583
      ("1000100101110011", '1', '1', "00", "111", "011", "001", '0', '-', "00"), -- i=2584
      ("1000100101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2585
      ("1001000101110011", '0', '1', "01", "111", "011", "001", '0', '-', "00"), -- i=2586
      ("1001100101110011", '1', '1', "01", "111", "011", "001", '0', '-', "00"), -- i=2587
      ("1001100101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2588
      ("1010000101110011", '0', '1', "10", "111", "011", "001", '0', '-', "00"), -- i=2589
      ("1010100101110011", '1', '1', "10", "111", "011", "001", '0', '-', "00"), -- i=2590
      ("1010100101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2591
      ("1011000101110011", '0', '1', "11", "111", "011", "001", '0', '-', "00"), -- i=2592
      ("1011100101110011", '1', '1', "11", "111", "011", "001", '0', '-', "00"), -- i=2593
      ("1011100101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2594
      ("0101000101110000", '0', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2595
      ("0101100101110000", '1', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2596
      ("0101100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2597
      ("0100000101110000", '0', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2598
      ("0100100101110000", '1', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2599
      ("0100100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2600
      ("0000000110011010", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2601
      ("0000100110011010", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2602
      ("0000100110011010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2603
      ("1000000101110100", '0', '1', "00", "111", "100", "001", '0', '-', "00"), -- i=2604
      ("1000100101110100", '1', '1', "00", "111", "100", "001", '0', '-', "00"), -- i=2605
      ("1000100101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2606
      ("1001000101110100", '0', '1', "01", "111", "100", "001", '0', '-', "00"), -- i=2607
      ("1001100101110100", '1', '1', "01", "111", "100", "001", '0', '-', "00"), -- i=2608
      ("1001100101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2609
      ("1010000101110100", '0', '1', "10", "111", "100", "001", '0', '-', "00"), -- i=2610
      ("1010100101110100", '1', '1', "10", "111", "100", "001", '0', '-', "00"), -- i=2611
      ("1010100101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2612
      ("1011000101110100", '0', '1', "11", "111", "100", "001", '0', '-', "00"), -- i=2613
      ("1011100101110100", '1', '1', "11", "111", "100", "001", '0', '-', "00"), -- i=2614
      ("1011100101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2615
      ("0101000101110000", '0', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2616
      ("0101100101110000", '1', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2617
      ("0101100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2618
      ("0100000101110000", '0', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2619
      ("0100100101110000", '1', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2620
      ("0100100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2621
      ("0000000100000100", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2622
      ("0000100100000100", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2623
      ("0000100100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2624
      ("1000000101110101", '0', '1', "00", "111", "101", "001", '0', '-', "00"), -- i=2625
      ("1000100101110101", '1', '1', "00", "111", "101", "001", '0', '-', "00"), -- i=2626
      ("1000100101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2627
      ("1001000101110101", '0', '1', "01", "111", "101", "001", '0', '-', "00"), -- i=2628
      ("1001100101110101", '1', '1', "01", "111", "101", "001", '0', '-', "00"), -- i=2629
      ("1001100101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2630
      ("1010000101110101", '0', '1', "10", "111", "101", "001", '0', '-', "00"), -- i=2631
      ("1010100101110101", '1', '1', "10", "111", "101", "001", '0', '-', "00"), -- i=2632
      ("1010100101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2633
      ("1011000101110101", '0', '1', "11", "111", "101", "001", '0', '-', "00"), -- i=2634
      ("1011100101110101", '1', '1', "11", "111", "101", "001", '0', '-', "00"), -- i=2635
      ("1011100101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2636
      ("0101000101110000", '0', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2637
      ("0101100101110000", '1', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2638
      ("0101100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2639
      ("0100000101110000", '0', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2640
      ("0100100101110000", '1', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2641
      ("0100100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2642
      ("0000000100110001", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2643
      ("0000100100110001", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2644
      ("0000100100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2645
      ("1000000101110110", '0', '1', "00", "111", "110", "001", '0', '-', "00"), -- i=2646
      ("1000100101110110", '1', '1', "00", "111", "110", "001", '0', '-', "00"), -- i=2647
      ("1000100101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2648
      ("1001000101110110", '0', '1', "01", "111", "110", "001", '0', '-', "00"), -- i=2649
      ("1001100101110110", '1', '1', "01", "111", "110", "001", '0', '-', "00"), -- i=2650
      ("1001100101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2651
      ("1010000101110110", '0', '1', "10", "111", "110", "001", '0', '-', "00"), -- i=2652
      ("1010100101110110", '1', '1', "10", "111", "110", "001", '0', '-', "00"), -- i=2653
      ("1010100101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2654
      ("1011000101110110", '0', '1', "11", "111", "110", "001", '0', '-', "00"), -- i=2655
      ("1011100101110110", '1', '1', "11", "111", "110", "001", '0', '-', "00"), -- i=2656
      ("1011100101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2657
      ("0101000101110000", '0', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2658
      ("0101100101110000", '1', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2659
      ("0101100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2660
      ("0100000101110000", '0', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2661
      ("0100100101110000", '1', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2662
      ("0100100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2663
      ("0000000110011100", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2664
      ("0000100110011100", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2665
      ("0000100110011100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2666
      ("1000000101110111", '0', '1', "00", "111", "111", "001", '0', '-', "00"), -- i=2667
      ("1000100101110111", '1', '1', "00", "111", "111", "001", '0', '-', "00"), -- i=2668
      ("1000100101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2669
      ("1001000101110111", '0', '1', "01", "111", "111", "001", '0', '-', "00"), -- i=2670
      ("1001100101110111", '1', '1', "01", "111", "111", "001", '0', '-', "00"), -- i=2671
      ("1001100101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2672
      ("1010000101110111", '0', '1', "10", "111", "111", "001", '0', '-', "00"), -- i=2673
      ("1010100101110111", '1', '1', "10", "111", "111", "001", '0', '-', "00"), -- i=2674
      ("1010100101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2675
      ("1011000101110111", '0', '1', "11", "111", "111", "001", '0', '-', "00"), -- i=2676
      ("1011100101110111", '1', '1', "11", "111", "111", "001", '0', '-', "00"), -- i=2677
      ("1011100101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2678
      ("0101000101110000", '0', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2679
      ("0101100101110000", '1', '1', "--", "111", "---", "001", '0', '1', "01"), -- i=2680
      ("0101100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2681
      ("0100000101110000", '0', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2682
      ("0100100101110000", '1', '0', "--", "111", "001", "---", '1', '-', "--"), -- i=2683
      ("0100100101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2684
      ("0000000101111110", '0', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2685
      ("0000100101111110", '1', '1', "--", "---", "---", "001", '0', '-', "10"), -- i=2686
      ("0000100101111110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2687
      ("1000001000000000", '0', '1', "00", "000", "000", "010", '0', '-', "00"), -- i=2688
      ("1000101000000000", '1', '1', "00", "000", "000", "010", '0', '-', "00"), -- i=2689
      ("1000101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2690
      ("1001001000000000", '0', '1', "01", "000", "000", "010", '0', '-', "00"), -- i=2691
      ("1001101000000000", '1', '1', "01", "000", "000", "010", '0', '-', "00"), -- i=2692
      ("1001101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2693
      ("1010001000000000", '0', '1', "10", "000", "000", "010", '0', '-', "00"), -- i=2694
      ("1010101000000000", '1', '1', "10", "000", "000", "010", '0', '-', "00"), -- i=2695
      ("1010101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2696
      ("1011001000000000", '0', '1', "11", "000", "000", "010", '0', '-', "00"), -- i=2697
      ("1011101000000000", '1', '1', "11", "000", "000", "010", '0', '-', "00"), -- i=2698
      ("1011101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2699
      ("0101001000000000", '0', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2700
      ("0101101000000000", '1', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2701
      ("0101101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2702
      ("0100001000000000", '0', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2703
      ("0100101000000000", '1', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2704
      ("0100101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2705
      ("0000001001110100", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2706
      ("0000101001110100", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2707
      ("0000101001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2708
      ("1000001000000001", '0', '1', "00", "000", "001", "010", '0', '-', "00"), -- i=2709
      ("1000101000000001", '1', '1', "00", "000", "001", "010", '0', '-', "00"), -- i=2710
      ("1000101000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2711
      ("1001001000000001", '0', '1', "01", "000", "001", "010", '0', '-', "00"), -- i=2712
      ("1001101000000001", '1', '1', "01", "000", "001", "010", '0', '-', "00"), -- i=2713
      ("1001101000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2714
      ("1010001000000001", '0', '1', "10", "000", "001", "010", '0', '-', "00"), -- i=2715
      ("1010101000000001", '1', '1', "10", "000", "001", "010", '0', '-', "00"), -- i=2716
      ("1010101000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2717
      ("1011001000000001", '0', '1', "11", "000", "001", "010", '0', '-', "00"), -- i=2718
      ("1011101000000001", '1', '1', "11", "000", "001", "010", '0', '-', "00"), -- i=2719
      ("1011101000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2720
      ("0101001000000000", '0', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2721
      ("0101101000000000", '1', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2722
      ("0101101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2723
      ("0100001000000000", '0', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2724
      ("0100101000000000", '1', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2725
      ("0100101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2726
      ("0000001001110001", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2727
      ("0000101001110001", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2728
      ("0000101001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2729
      ("1000001000000010", '0', '1', "00", "000", "010", "010", '0', '-', "00"), -- i=2730
      ("1000101000000010", '1', '1', "00", "000", "010", "010", '0', '-', "00"), -- i=2731
      ("1000101000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2732
      ("1001001000000010", '0', '1', "01", "000", "010", "010", '0', '-', "00"), -- i=2733
      ("1001101000000010", '1', '1', "01", "000", "010", "010", '0', '-', "00"), -- i=2734
      ("1001101000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2735
      ("1010001000000010", '0', '1', "10", "000", "010", "010", '0', '-', "00"), -- i=2736
      ("1010101000000010", '1', '1', "10", "000", "010", "010", '0', '-', "00"), -- i=2737
      ("1010101000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2738
      ("1011001000000010", '0', '1', "11", "000", "010", "010", '0', '-', "00"), -- i=2739
      ("1011101000000010", '1', '1', "11", "000", "010", "010", '0', '-', "00"), -- i=2740
      ("1011101000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2741
      ("0101001000000000", '0', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2742
      ("0101101000000000", '1', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2743
      ("0101101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2744
      ("0100001000000000", '0', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2745
      ("0100101000000000", '1', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2746
      ("0100101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2747
      ("0000001010110000", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2748
      ("0000101010110000", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2749
      ("0000101010110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2750
      ("1000001000000011", '0', '1', "00", "000", "011", "010", '0', '-', "00"), -- i=2751
      ("1000101000000011", '1', '1', "00", "000", "011", "010", '0', '-', "00"), -- i=2752
      ("1000101000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2753
      ("1001001000000011", '0', '1', "01", "000", "011", "010", '0', '-', "00"), -- i=2754
      ("1001101000000011", '1', '1', "01", "000", "011", "010", '0', '-', "00"), -- i=2755
      ("1001101000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2756
      ("1010001000000011", '0', '1', "10", "000", "011", "010", '0', '-', "00"), -- i=2757
      ("1010101000000011", '1', '1', "10", "000", "011", "010", '0', '-', "00"), -- i=2758
      ("1010101000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2759
      ("1011001000000011", '0', '1', "11", "000", "011", "010", '0', '-', "00"), -- i=2760
      ("1011101000000011", '1', '1', "11", "000", "011", "010", '0', '-', "00"), -- i=2761
      ("1011101000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2762
      ("0101001000000000", '0', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2763
      ("0101101000000000", '1', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2764
      ("0101101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2765
      ("0100001000000000", '0', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2766
      ("0100101000000000", '1', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2767
      ("0100101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2768
      ("0000001010000000", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2769
      ("0000101010000000", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2770
      ("0000101010000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2771
      ("1000001000000100", '0', '1', "00", "000", "100", "010", '0', '-', "00"), -- i=2772
      ("1000101000000100", '1', '1', "00", "000", "100", "010", '0', '-', "00"), -- i=2773
      ("1000101000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2774
      ("1001001000000100", '0', '1', "01", "000", "100", "010", '0', '-', "00"), -- i=2775
      ("1001101000000100", '1', '1', "01", "000", "100", "010", '0', '-', "00"), -- i=2776
      ("1001101000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2777
      ("1010001000000100", '0', '1', "10", "000", "100", "010", '0', '-', "00"), -- i=2778
      ("1010101000000100", '1', '1', "10", "000", "100", "010", '0', '-', "00"), -- i=2779
      ("1010101000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2780
      ("1011001000000100", '0', '1', "11", "000", "100", "010", '0', '-', "00"), -- i=2781
      ("1011101000000100", '1', '1', "11", "000", "100", "010", '0', '-', "00"), -- i=2782
      ("1011101000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2783
      ("0101001000000000", '0', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2784
      ("0101101000000000", '1', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2785
      ("0101101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2786
      ("0100001000000000", '0', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2787
      ("0100101000000000", '1', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2788
      ("0100101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2789
      ("0000001000000110", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2790
      ("0000101000000110", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2791
      ("0000101000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2792
      ("1000001000000101", '0', '1', "00", "000", "101", "010", '0', '-', "00"), -- i=2793
      ("1000101000000101", '1', '1', "00", "000", "101", "010", '0', '-', "00"), -- i=2794
      ("1000101000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2795
      ("1001001000000101", '0', '1', "01", "000", "101", "010", '0', '-', "00"), -- i=2796
      ("1001101000000101", '1', '1', "01", "000", "101", "010", '0', '-', "00"), -- i=2797
      ("1001101000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2798
      ("1010001000000101", '0', '1', "10", "000", "101", "010", '0', '-', "00"), -- i=2799
      ("1010101000000101", '1', '1', "10", "000", "101", "010", '0', '-', "00"), -- i=2800
      ("1010101000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2801
      ("1011001000000101", '0', '1', "11", "000", "101", "010", '0', '-', "00"), -- i=2802
      ("1011101000000101", '1', '1', "11", "000", "101", "010", '0', '-', "00"), -- i=2803
      ("1011101000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2804
      ("0101001000000000", '0', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2805
      ("0101101000000000", '1', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2806
      ("0101101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2807
      ("0100001000000000", '0', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2808
      ("0100101000000000", '1', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2809
      ("0100101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2810
      ("0000001000001111", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2811
      ("0000101000001111", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2812
      ("0000101000001111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2813
      ("1000001000000110", '0', '1', "00", "000", "110", "010", '0', '-', "00"), -- i=2814
      ("1000101000000110", '1', '1', "00", "000", "110", "010", '0', '-', "00"), -- i=2815
      ("1000101000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2816
      ("1001001000000110", '0', '1', "01", "000", "110", "010", '0', '-', "00"), -- i=2817
      ("1001101000000110", '1', '1', "01", "000", "110", "010", '0', '-', "00"), -- i=2818
      ("1001101000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2819
      ("1010001000000110", '0', '1', "10", "000", "110", "010", '0', '-', "00"), -- i=2820
      ("1010101000000110", '1', '1', "10", "000", "110", "010", '0', '-', "00"), -- i=2821
      ("1010101000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2822
      ("1011001000000110", '0', '1', "11", "000", "110", "010", '0', '-', "00"), -- i=2823
      ("1011101000000110", '1', '1', "11", "000", "110", "010", '0', '-', "00"), -- i=2824
      ("1011101000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2825
      ("0101001000000000", '0', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2826
      ("0101101000000000", '1', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2827
      ("0101101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2828
      ("0100001000000000", '0', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2829
      ("0100101000000000", '1', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2830
      ("0100101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2831
      ("0000001010100011", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2832
      ("0000101010100011", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2833
      ("0000101010100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2834
      ("1000001000000111", '0', '1', "00", "000", "111", "010", '0', '-', "00"), -- i=2835
      ("1000101000000111", '1', '1', "00", "000", "111", "010", '0', '-', "00"), -- i=2836
      ("1000101000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2837
      ("1001001000000111", '0', '1', "01", "000", "111", "010", '0', '-', "00"), -- i=2838
      ("1001101000000111", '1', '1', "01", "000", "111", "010", '0', '-', "00"), -- i=2839
      ("1001101000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2840
      ("1010001000000111", '0', '1', "10", "000", "111", "010", '0', '-', "00"), -- i=2841
      ("1010101000000111", '1', '1', "10", "000", "111", "010", '0', '-', "00"), -- i=2842
      ("1010101000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2843
      ("1011001000000111", '0', '1', "11", "000", "111", "010", '0', '-', "00"), -- i=2844
      ("1011101000000111", '1', '1', "11", "000", "111", "010", '0', '-', "00"), -- i=2845
      ("1011101000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2846
      ("0101001000000000", '0', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2847
      ("0101101000000000", '1', '1', "--", "000", "---", "010", '0', '1', "01"), -- i=2848
      ("0101101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2849
      ("0100001000000000", '0', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2850
      ("0100101000000000", '1', '0', "--", "000", "010", "---", '1', '-', "--"), -- i=2851
      ("0100101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2852
      ("0000001000001101", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2853
      ("0000101000001101", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2854
      ("0000101000001101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2855
      ("1000001000010000", '0', '1', "00", "001", "000", "010", '0', '-', "00"), -- i=2856
      ("1000101000010000", '1', '1', "00", "001", "000", "010", '0', '-', "00"), -- i=2857
      ("1000101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2858
      ("1001001000010000", '0', '1', "01", "001", "000", "010", '0', '-', "00"), -- i=2859
      ("1001101000010000", '1', '1', "01", "001", "000", "010", '0', '-', "00"), -- i=2860
      ("1001101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2861
      ("1010001000010000", '0', '1', "10", "001", "000", "010", '0', '-', "00"), -- i=2862
      ("1010101000010000", '1', '1', "10", "001", "000", "010", '0', '-', "00"), -- i=2863
      ("1010101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2864
      ("1011001000010000", '0', '1', "11", "001", "000", "010", '0', '-', "00"), -- i=2865
      ("1011101000010000", '1', '1', "11", "001", "000", "010", '0', '-', "00"), -- i=2866
      ("1011101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2867
      ("0101001000010000", '0', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=2868
      ("0101101000010000", '1', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=2869
      ("0101101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2870
      ("0100001000010000", '0', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=2871
      ("0100101000010000", '1', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=2872
      ("0100101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2873
      ("0000001011001110", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2874
      ("0000101011001110", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2875
      ("0000101011001110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2876
      ("1000001000010001", '0', '1', "00", "001", "001", "010", '0', '-', "00"), -- i=2877
      ("1000101000010001", '1', '1', "00", "001", "001", "010", '0', '-', "00"), -- i=2878
      ("1000101000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2879
      ("1001001000010001", '0', '1', "01", "001", "001", "010", '0', '-', "00"), -- i=2880
      ("1001101000010001", '1', '1', "01", "001", "001", "010", '0', '-', "00"), -- i=2881
      ("1001101000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2882
      ("1010001000010001", '0', '1', "10", "001", "001", "010", '0', '-', "00"), -- i=2883
      ("1010101000010001", '1', '1', "10", "001", "001", "010", '0', '-', "00"), -- i=2884
      ("1010101000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2885
      ("1011001000010001", '0', '1', "11", "001", "001", "010", '0', '-', "00"), -- i=2886
      ("1011101000010001", '1', '1', "11", "001", "001", "010", '0', '-', "00"), -- i=2887
      ("1011101000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2888
      ("0101001000010000", '0', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=2889
      ("0101101000010000", '1', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=2890
      ("0101101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2891
      ("0100001000010000", '0', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=2892
      ("0100101000010000", '1', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=2893
      ("0100101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2894
      ("0000001010101100", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2895
      ("0000101010101100", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2896
      ("0000101010101100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2897
      ("1000001000010010", '0', '1', "00", "001", "010", "010", '0', '-', "00"), -- i=2898
      ("1000101000010010", '1', '1', "00", "001", "010", "010", '0', '-', "00"), -- i=2899
      ("1000101000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2900
      ("1001001000010010", '0', '1', "01", "001", "010", "010", '0', '-', "00"), -- i=2901
      ("1001101000010010", '1', '1', "01", "001", "010", "010", '0', '-', "00"), -- i=2902
      ("1001101000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2903
      ("1010001000010010", '0', '1', "10", "001", "010", "010", '0', '-', "00"), -- i=2904
      ("1010101000010010", '1', '1', "10", "001", "010", "010", '0', '-', "00"), -- i=2905
      ("1010101000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2906
      ("1011001000010010", '0', '1', "11", "001", "010", "010", '0', '-', "00"), -- i=2907
      ("1011101000010010", '1', '1', "11", "001", "010", "010", '0', '-', "00"), -- i=2908
      ("1011101000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2909
      ("0101001000010000", '0', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=2910
      ("0101101000010000", '1', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=2911
      ("0101101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2912
      ("0100001000010000", '0', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=2913
      ("0100101000010000", '1', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=2914
      ("0100101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2915
      ("0000001011100101", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2916
      ("0000101011100101", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2917
      ("0000101011100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2918
      ("1000001000010011", '0', '1', "00", "001", "011", "010", '0', '-', "00"), -- i=2919
      ("1000101000010011", '1', '1', "00", "001", "011", "010", '0', '-', "00"), -- i=2920
      ("1000101000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2921
      ("1001001000010011", '0', '1', "01", "001", "011", "010", '0', '-', "00"), -- i=2922
      ("1001101000010011", '1', '1', "01", "001", "011", "010", '0', '-', "00"), -- i=2923
      ("1001101000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2924
      ("1010001000010011", '0', '1', "10", "001", "011", "010", '0', '-', "00"), -- i=2925
      ("1010101000010011", '1', '1', "10", "001", "011", "010", '0', '-', "00"), -- i=2926
      ("1010101000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2927
      ("1011001000010011", '0', '1', "11", "001", "011", "010", '0', '-', "00"), -- i=2928
      ("1011101000010011", '1', '1', "11", "001", "011", "010", '0', '-', "00"), -- i=2929
      ("1011101000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2930
      ("0101001000010000", '0', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=2931
      ("0101101000010000", '1', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=2932
      ("0101101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2933
      ("0100001000010000", '0', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=2934
      ("0100101000010000", '1', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=2935
      ("0100101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2936
      ("0000001001111100", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2937
      ("0000101001111100", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2938
      ("0000101001111100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2939
      ("1000001000010100", '0', '1', "00", "001", "100", "010", '0', '-', "00"), -- i=2940
      ("1000101000010100", '1', '1', "00", "001", "100", "010", '0', '-', "00"), -- i=2941
      ("1000101000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2942
      ("1001001000010100", '0', '1', "01", "001", "100", "010", '0', '-', "00"), -- i=2943
      ("1001101000010100", '1', '1', "01", "001", "100", "010", '0', '-', "00"), -- i=2944
      ("1001101000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2945
      ("1010001000010100", '0', '1', "10", "001", "100", "010", '0', '-', "00"), -- i=2946
      ("1010101000010100", '1', '1', "10", "001", "100", "010", '0', '-', "00"), -- i=2947
      ("1010101000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2948
      ("1011001000010100", '0', '1', "11", "001", "100", "010", '0', '-', "00"), -- i=2949
      ("1011101000010100", '1', '1', "11", "001", "100", "010", '0', '-', "00"), -- i=2950
      ("1011101000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2951
      ("0101001000010000", '0', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=2952
      ("0101101000010000", '1', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=2953
      ("0101101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2954
      ("0100001000010000", '0', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=2955
      ("0100101000010000", '1', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=2956
      ("0100101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2957
      ("0000001000000000", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2958
      ("0000101000000000", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2959
      ("0000101000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2960
      ("1000001000010101", '0', '1', "00", "001", "101", "010", '0', '-', "00"), -- i=2961
      ("1000101000010101", '1', '1', "00", "001", "101", "010", '0', '-', "00"), -- i=2962
      ("1000101000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2963
      ("1001001000010101", '0', '1', "01", "001", "101", "010", '0', '-', "00"), -- i=2964
      ("1001101000010101", '1', '1', "01", "001", "101", "010", '0', '-', "00"), -- i=2965
      ("1001101000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2966
      ("1010001000010101", '0', '1', "10", "001", "101", "010", '0', '-', "00"), -- i=2967
      ("1010101000010101", '1', '1', "10", "001", "101", "010", '0', '-', "00"), -- i=2968
      ("1010101000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2969
      ("1011001000010101", '0', '1', "11", "001", "101", "010", '0', '-', "00"), -- i=2970
      ("1011101000010101", '1', '1', "11", "001", "101", "010", '0', '-', "00"), -- i=2971
      ("1011101000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2972
      ("0101001000010000", '0', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=2973
      ("0101101000010000", '1', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=2974
      ("0101101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2975
      ("0100001000010000", '0', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=2976
      ("0100101000010000", '1', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=2977
      ("0100101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2978
      ("0000001011101001", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2979
      ("0000101011101001", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=2980
      ("0000101011101001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2981
      ("1000001000010110", '0', '1', "00", "001", "110", "010", '0', '-', "00"), -- i=2982
      ("1000101000010110", '1', '1', "00", "001", "110", "010", '0', '-', "00"), -- i=2983
      ("1000101000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2984
      ("1001001000010110", '0', '1', "01", "001", "110", "010", '0', '-', "00"), -- i=2985
      ("1001101000010110", '1', '1', "01", "001", "110", "010", '0', '-', "00"), -- i=2986
      ("1001101000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2987
      ("1010001000010110", '0', '1', "10", "001", "110", "010", '0', '-', "00"), -- i=2988
      ("1010101000010110", '1', '1', "10", "001", "110", "010", '0', '-', "00"), -- i=2989
      ("1010101000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2990
      ("1011001000010110", '0', '1', "11", "001", "110", "010", '0', '-', "00"), -- i=2991
      ("1011101000010110", '1', '1', "11", "001", "110", "010", '0', '-', "00"), -- i=2992
      ("1011101000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2993
      ("0101001000010000", '0', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=2994
      ("0101101000010000", '1', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=2995
      ("0101101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2996
      ("0100001000010000", '0', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=2997
      ("0100101000010000", '1', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=2998
      ("0100101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=2999
      ("0000001010000001", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3000
      ("0000101010000001", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3001
      ("0000101010000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3002
      ("1000001000010111", '0', '1', "00", "001", "111", "010", '0', '-', "00"), -- i=3003
      ("1000101000010111", '1', '1', "00", "001", "111", "010", '0', '-', "00"), -- i=3004
      ("1000101000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3005
      ("1001001000010111", '0', '1', "01", "001", "111", "010", '0', '-', "00"), -- i=3006
      ("1001101000010111", '1', '1', "01", "001", "111", "010", '0', '-', "00"), -- i=3007
      ("1001101000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3008
      ("1010001000010111", '0', '1', "10", "001", "111", "010", '0', '-', "00"), -- i=3009
      ("1010101000010111", '1', '1', "10", "001", "111", "010", '0', '-', "00"), -- i=3010
      ("1010101000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3011
      ("1011001000010111", '0', '1', "11", "001", "111", "010", '0', '-', "00"), -- i=3012
      ("1011101000010111", '1', '1', "11", "001", "111", "010", '0', '-', "00"), -- i=3013
      ("1011101000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3014
      ("0101001000010000", '0', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=3015
      ("0101101000010000", '1', '1', "--", "001", "---", "010", '0', '1', "01"), -- i=3016
      ("0101101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3017
      ("0100001000010000", '0', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=3018
      ("0100101000010000", '1', '0', "--", "001", "010", "---", '1', '-', "--"), -- i=3019
      ("0100101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3020
      ("0000001011011111", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3021
      ("0000101011011111", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3022
      ("0000101011011111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3023
      ("1000001000100000", '0', '1', "00", "010", "000", "010", '0', '-', "00"), -- i=3024
      ("1000101000100000", '1', '1', "00", "010", "000", "010", '0', '-', "00"), -- i=3025
      ("1000101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3026
      ("1001001000100000", '0', '1', "01", "010", "000", "010", '0', '-', "00"), -- i=3027
      ("1001101000100000", '1', '1', "01", "010", "000", "010", '0', '-', "00"), -- i=3028
      ("1001101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3029
      ("1010001000100000", '0', '1', "10", "010", "000", "010", '0', '-', "00"), -- i=3030
      ("1010101000100000", '1', '1', "10", "010", "000", "010", '0', '-', "00"), -- i=3031
      ("1010101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3032
      ("1011001000100000", '0', '1', "11", "010", "000", "010", '0', '-', "00"), -- i=3033
      ("1011101000100000", '1', '1', "11", "010", "000", "010", '0', '-', "00"), -- i=3034
      ("1011101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3035
      ("0101001000100000", '0', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3036
      ("0101101000100000", '1', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3037
      ("0101101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3038
      ("0100001000100000", '0', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3039
      ("0100101000100000", '1', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3040
      ("0100101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3041
      ("0000001010101111", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3042
      ("0000101010101111", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3043
      ("0000101010101111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3044
      ("1000001000100001", '0', '1', "00", "010", "001", "010", '0', '-', "00"), -- i=3045
      ("1000101000100001", '1', '1', "00", "010", "001", "010", '0', '-', "00"), -- i=3046
      ("1000101000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3047
      ("1001001000100001", '0', '1', "01", "010", "001", "010", '0', '-', "00"), -- i=3048
      ("1001101000100001", '1', '1', "01", "010", "001", "010", '0', '-', "00"), -- i=3049
      ("1001101000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3050
      ("1010001000100001", '0', '1', "10", "010", "001", "010", '0', '-', "00"), -- i=3051
      ("1010101000100001", '1', '1', "10", "010", "001", "010", '0', '-', "00"), -- i=3052
      ("1010101000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3053
      ("1011001000100001", '0', '1', "11", "010", "001", "010", '0', '-', "00"), -- i=3054
      ("1011101000100001", '1', '1', "11", "010", "001", "010", '0', '-', "00"), -- i=3055
      ("1011101000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3056
      ("0101001000100000", '0', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3057
      ("0101101000100000", '1', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3058
      ("0101101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3059
      ("0100001000100000", '0', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3060
      ("0100101000100000", '1', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3061
      ("0100101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3062
      ("0000001001010100", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3063
      ("0000101001010100", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3064
      ("0000101001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3065
      ("1000001000100010", '0', '1', "00", "010", "010", "010", '0', '-', "00"), -- i=3066
      ("1000101000100010", '1', '1', "00", "010", "010", "010", '0', '-', "00"), -- i=3067
      ("1000101000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3068
      ("1001001000100010", '0', '1', "01", "010", "010", "010", '0', '-', "00"), -- i=3069
      ("1001101000100010", '1', '1', "01", "010", "010", "010", '0', '-', "00"), -- i=3070
      ("1001101000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3071
      ("1010001000100010", '0', '1', "10", "010", "010", "010", '0', '-', "00"), -- i=3072
      ("1010101000100010", '1', '1', "10", "010", "010", "010", '0', '-', "00"), -- i=3073
      ("1010101000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3074
      ("1011001000100010", '0', '1', "11", "010", "010", "010", '0', '-', "00"), -- i=3075
      ("1011101000100010", '1', '1', "11", "010", "010", "010", '0', '-', "00"), -- i=3076
      ("1011101000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3077
      ("0101001000100000", '0', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3078
      ("0101101000100000", '1', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3079
      ("0101101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3080
      ("0100001000100000", '0', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3081
      ("0100101000100000", '1', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3082
      ("0100101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3083
      ("0000001001000110", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3084
      ("0000101001000110", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3085
      ("0000101001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3086
      ("1000001000100011", '0', '1', "00", "010", "011", "010", '0', '-', "00"), -- i=3087
      ("1000101000100011", '1', '1', "00", "010", "011", "010", '0', '-', "00"), -- i=3088
      ("1000101000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3089
      ("1001001000100011", '0', '1', "01", "010", "011", "010", '0', '-', "00"), -- i=3090
      ("1001101000100011", '1', '1', "01", "010", "011", "010", '0', '-', "00"), -- i=3091
      ("1001101000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3092
      ("1010001000100011", '0', '1', "10", "010", "011", "010", '0', '-', "00"), -- i=3093
      ("1010101000100011", '1', '1', "10", "010", "011", "010", '0', '-', "00"), -- i=3094
      ("1010101000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3095
      ("1011001000100011", '0', '1', "11", "010", "011", "010", '0', '-', "00"), -- i=3096
      ("1011101000100011", '1', '1', "11", "010", "011", "010", '0', '-', "00"), -- i=3097
      ("1011101000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3098
      ("0101001000100000", '0', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3099
      ("0101101000100000", '1', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3100
      ("0101101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3101
      ("0100001000100000", '0', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3102
      ("0100101000100000", '1', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3103
      ("0100101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3104
      ("0000001000100110", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3105
      ("0000101000100110", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3106
      ("0000101000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3107
      ("1000001000100100", '0', '1', "00", "010", "100", "010", '0', '-', "00"), -- i=3108
      ("1000101000100100", '1', '1', "00", "010", "100", "010", '0', '-', "00"), -- i=3109
      ("1000101000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3110
      ("1001001000100100", '0', '1', "01", "010", "100", "010", '0', '-', "00"), -- i=3111
      ("1001101000100100", '1', '1', "01", "010", "100", "010", '0', '-', "00"), -- i=3112
      ("1001101000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3113
      ("1010001000100100", '0', '1', "10", "010", "100", "010", '0', '-', "00"), -- i=3114
      ("1010101000100100", '1', '1', "10", "010", "100", "010", '0', '-', "00"), -- i=3115
      ("1010101000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3116
      ("1011001000100100", '0', '1', "11", "010", "100", "010", '0', '-', "00"), -- i=3117
      ("1011101000100100", '1', '1', "11", "010", "100", "010", '0', '-', "00"), -- i=3118
      ("1011101000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3119
      ("0101001000100000", '0', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3120
      ("0101101000100000", '1', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3121
      ("0101101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3122
      ("0100001000100000", '0', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3123
      ("0100101000100000", '1', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3124
      ("0100101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3125
      ("0000001010101001", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3126
      ("0000101010101001", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3127
      ("0000101010101001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3128
      ("1000001000100101", '0', '1', "00", "010", "101", "010", '0', '-', "00"), -- i=3129
      ("1000101000100101", '1', '1', "00", "010", "101", "010", '0', '-', "00"), -- i=3130
      ("1000101000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3131
      ("1001001000100101", '0', '1', "01", "010", "101", "010", '0', '-', "00"), -- i=3132
      ("1001101000100101", '1', '1', "01", "010", "101", "010", '0', '-', "00"), -- i=3133
      ("1001101000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3134
      ("1010001000100101", '0', '1', "10", "010", "101", "010", '0', '-', "00"), -- i=3135
      ("1010101000100101", '1', '1', "10", "010", "101", "010", '0', '-', "00"), -- i=3136
      ("1010101000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3137
      ("1011001000100101", '0', '1', "11", "010", "101", "010", '0', '-', "00"), -- i=3138
      ("1011101000100101", '1', '1', "11", "010", "101", "010", '0', '-', "00"), -- i=3139
      ("1011101000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3140
      ("0101001000100000", '0', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3141
      ("0101101000100000", '1', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3142
      ("0101101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3143
      ("0100001000100000", '0', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3144
      ("0100101000100000", '1', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3145
      ("0100101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3146
      ("0000001011111010", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3147
      ("0000101011111010", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3148
      ("0000101011111010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3149
      ("1000001000100110", '0', '1', "00", "010", "110", "010", '0', '-', "00"), -- i=3150
      ("1000101000100110", '1', '1', "00", "010", "110", "010", '0', '-', "00"), -- i=3151
      ("1000101000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3152
      ("1001001000100110", '0', '1', "01", "010", "110", "010", '0', '-', "00"), -- i=3153
      ("1001101000100110", '1', '1', "01", "010", "110", "010", '0', '-', "00"), -- i=3154
      ("1001101000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3155
      ("1010001000100110", '0', '1', "10", "010", "110", "010", '0', '-', "00"), -- i=3156
      ("1010101000100110", '1', '1', "10", "010", "110", "010", '0', '-', "00"), -- i=3157
      ("1010101000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3158
      ("1011001000100110", '0', '1', "11", "010", "110", "010", '0', '-', "00"), -- i=3159
      ("1011101000100110", '1', '1', "11", "010", "110", "010", '0', '-', "00"), -- i=3160
      ("1011101000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3161
      ("0101001000100000", '0', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3162
      ("0101101000100000", '1', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3163
      ("0101101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3164
      ("0100001000100000", '0', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3165
      ("0100101000100000", '1', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3166
      ("0100101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3167
      ("0000001010101001", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3168
      ("0000101010101001", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3169
      ("0000101010101001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3170
      ("1000001000100111", '0', '1', "00", "010", "111", "010", '0', '-', "00"), -- i=3171
      ("1000101000100111", '1', '1', "00", "010", "111", "010", '0', '-', "00"), -- i=3172
      ("1000101000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3173
      ("1001001000100111", '0', '1', "01", "010", "111", "010", '0', '-', "00"), -- i=3174
      ("1001101000100111", '1', '1', "01", "010", "111", "010", '0', '-', "00"), -- i=3175
      ("1001101000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3176
      ("1010001000100111", '0', '1', "10", "010", "111", "010", '0', '-', "00"), -- i=3177
      ("1010101000100111", '1', '1', "10", "010", "111", "010", '0', '-', "00"), -- i=3178
      ("1010101000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3179
      ("1011001000100111", '0', '1', "11", "010", "111", "010", '0', '-', "00"), -- i=3180
      ("1011101000100111", '1', '1', "11", "010", "111", "010", '0', '-', "00"), -- i=3181
      ("1011101000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3182
      ("0101001000100000", '0', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3183
      ("0101101000100000", '1', '1', "--", "010", "---", "010", '0', '1', "01"), -- i=3184
      ("0101101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3185
      ("0100001000100000", '0', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3186
      ("0100101000100000", '1', '0', "--", "010", "010", "---", '1', '-', "--"), -- i=3187
      ("0100101000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3188
      ("0000001000000010", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3189
      ("0000101000000010", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3190
      ("0000101000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3191
      ("1000001000110000", '0', '1', "00", "011", "000", "010", '0', '-', "00"), -- i=3192
      ("1000101000110000", '1', '1', "00", "011", "000", "010", '0', '-', "00"), -- i=3193
      ("1000101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3194
      ("1001001000110000", '0', '1', "01", "011", "000", "010", '0', '-', "00"), -- i=3195
      ("1001101000110000", '1', '1', "01", "011", "000", "010", '0', '-', "00"), -- i=3196
      ("1001101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3197
      ("1010001000110000", '0', '1', "10", "011", "000", "010", '0', '-', "00"), -- i=3198
      ("1010101000110000", '1', '1', "10", "011", "000", "010", '0', '-', "00"), -- i=3199
      ("1010101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3200
      ("1011001000110000", '0', '1', "11", "011", "000", "010", '0', '-', "00"), -- i=3201
      ("1011101000110000", '1', '1', "11", "011", "000", "010", '0', '-', "00"), -- i=3202
      ("1011101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3203
      ("0101001000110000", '0', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3204
      ("0101101000110000", '1', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3205
      ("0101101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3206
      ("0100001000110000", '0', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3207
      ("0100101000110000", '1', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3208
      ("0100101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3209
      ("0000001000011011", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3210
      ("0000101000011011", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3211
      ("0000101000011011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3212
      ("1000001000110001", '0', '1', "00", "011", "001", "010", '0', '-', "00"), -- i=3213
      ("1000101000110001", '1', '1', "00", "011", "001", "010", '0', '-', "00"), -- i=3214
      ("1000101000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3215
      ("1001001000110001", '0', '1', "01", "011", "001", "010", '0', '-', "00"), -- i=3216
      ("1001101000110001", '1', '1', "01", "011", "001", "010", '0', '-', "00"), -- i=3217
      ("1001101000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3218
      ("1010001000110001", '0', '1', "10", "011", "001", "010", '0', '-', "00"), -- i=3219
      ("1010101000110001", '1', '1', "10", "011", "001", "010", '0', '-', "00"), -- i=3220
      ("1010101000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3221
      ("1011001000110001", '0', '1', "11", "011", "001", "010", '0', '-', "00"), -- i=3222
      ("1011101000110001", '1', '1', "11", "011", "001", "010", '0', '-', "00"), -- i=3223
      ("1011101000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3224
      ("0101001000110000", '0', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3225
      ("0101101000110000", '1', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3226
      ("0101101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3227
      ("0100001000110000", '0', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3228
      ("0100101000110000", '1', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3229
      ("0100101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3230
      ("0000001001000001", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3231
      ("0000101001000001", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3232
      ("0000101001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3233
      ("1000001000110010", '0', '1', "00", "011", "010", "010", '0', '-', "00"), -- i=3234
      ("1000101000110010", '1', '1', "00", "011", "010", "010", '0', '-', "00"), -- i=3235
      ("1000101000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3236
      ("1001001000110010", '0', '1', "01", "011", "010", "010", '0', '-', "00"), -- i=3237
      ("1001101000110010", '1', '1', "01", "011", "010", "010", '0', '-', "00"), -- i=3238
      ("1001101000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3239
      ("1010001000110010", '0', '1', "10", "011", "010", "010", '0', '-', "00"), -- i=3240
      ("1010101000110010", '1', '1', "10", "011", "010", "010", '0', '-', "00"), -- i=3241
      ("1010101000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3242
      ("1011001000110010", '0', '1', "11", "011", "010", "010", '0', '-', "00"), -- i=3243
      ("1011101000110010", '1', '1', "11", "011", "010", "010", '0', '-', "00"), -- i=3244
      ("1011101000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3245
      ("0101001000110000", '0', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3246
      ("0101101000110000", '1', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3247
      ("0101101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3248
      ("0100001000110000", '0', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3249
      ("0100101000110000", '1', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3250
      ("0100101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3251
      ("0000001001000001", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3252
      ("0000101001000001", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3253
      ("0000101001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3254
      ("1000001000110011", '0', '1', "00", "011", "011", "010", '0', '-', "00"), -- i=3255
      ("1000101000110011", '1', '1', "00", "011", "011", "010", '0', '-', "00"), -- i=3256
      ("1000101000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3257
      ("1001001000110011", '0', '1', "01", "011", "011", "010", '0', '-', "00"), -- i=3258
      ("1001101000110011", '1', '1', "01", "011", "011", "010", '0', '-', "00"), -- i=3259
      ("1001101000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3260
      ("1010001000110011", '0', '1', "10", "011", "011", "010", '0', '-', "00"), -- i=3261
      ("1010101000110011", '1', '1', "10", "011", "011", "010", '0', '-', "00"), -- i=3262
      ("1010101000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3263
      ("1011001000110011", '0', '1', "11", "011", "011", "010", '0', '-', "00"), -- i=3264
      ("1011101000110011", '1', '1', "11", "011", "011", "010", '0', '-', "00"), -- i=3265
      ("1011101000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3266
      ("0101001000110000", '0', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3267
      ("0101101000110000", '1', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3268
      ("0101101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3269
      ("0100001000110000", '0', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3270
      ("0100101000110000", '1', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3271
      ("0100101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3272
      ("0000001001010000", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3273
      ("0000101001010000", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3274
      ("0000101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3275
      ("1000001000110100", '0', '1', "00", "011", "100", "010", '0', '-', "00"), -- i=3276
      ("1000101000110100", '1', '1', "00", "011", "100", "010", '0', '-', "00"), -- i=3277
      ("1000101000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3278
      ("1001001000110100", '0', '1', "01", "011", "100", "010", '0', '-', "00"), -- i=3279
      ("1001101000110100", '1', '1', "01", "011", "100", "010", '0', '-', "00"), -- i=3280
      ("1001101000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3281
      ("1010001000110100", '0', '1', "10", "011", "100", "010", '0', '-', "00"), -- i=3282
      ("1010101000110100", '1', '1', "10", "011", "100", "010", '0', '-', "00"), -- i=3283
      ("1010101000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3284
      ("1011001000110100", '0', '1', "11", "011", "100", "010", '0', '-', "00"), -- i=3285
      ("1011101000110100", '1', '1', "11", "011", "100", "010", '0', '-', "00"), -- i=3286
      ("1011101000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3287
      ("0101001000110000", '0', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3288
      ("0101101000110000", '1', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3289
      ("0101101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3290
      ("0100001000110000", '0', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3291
      ("0100101000110000", '1', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3292
      ("0100101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3293
      ("0000001010100011", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3294
      ("0000101010100011", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3295
      ("0000101010100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3296
      ("1000001000110101", '0', '1', "00", "011", "101", "010", '0', '-', "00"), -- i=3297
      ("1000101000110101", '1', '1', "00", "011", "101", "010", '0', '-', "00"), -- i=3298
      ("1000101000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3299
      ("1001001000110101", '0', '1', "01", "011", "101", "010", '0', '-', "00"), -- i=3300
      ("1001101000110101", '1', '1', "01", "011", "101", "010", '0', '-', "00"), -- i=3301
      ("1001101000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3302
      ("1010001000110101", '0', '1', "10", "011", "101", "010", '0', '-', "00"), -- i=3303
      ("1010101000110101", '1', '1', "10", "011", "101", "010", '0', '-', "00"), -- i=3304
      ("1010101000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3305
      ("1011001000110101", '0', '1', "11", "011", "101", "010", '0', '-', "00"), -- i=3306
      ("1011101000110101", '1', '1', "11", "011", "101", "010", '0', '-', "00"), -- i=3307
      ("1011101000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3308
      ("0101001000110000", '0', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3309
      ("0101101000110000", '1', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3310
      ("0101101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3311
      ("0100001000110000", '0', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3312
      ("0100101000110000", '1', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3313
      ("0100101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3314
      ("0000001000011010", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3315
      ("0000101000011010", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3316
      ("0000101000011010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3317
      ("1000001000110110", '0', '1', "00", "011", "110", "010", '0', '-', "00"), -- i=3318
      ("1000101000110110", '1', '1', "00", "011", "110", "010", '0', '-', "00"), -- i=3319
      ("1000101000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3320
      ("1001001000110110", '0', '1', "01", "011", "110", "010", '0', '-', "00"), -- i=3321
      ("1001101000110110", '1', '1', "01", "011", "110", "010", '0', '-', "00"), -- i=3322
      ("1001101000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3323
      ("1010001000110110", '0', '1', "10", "011", "110", "010", '0', '-', "00"), -- i=3324
      ("1010101000110110", '1', '1', "10", "011", "110", "010", '0', '-', "00"), -- i=3325
      ("1010101000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3326
      ("1011001000110110", '0', '1', "11", "011", "110", "010", '0', '-', "00"), -- i=3327
      ("1011101000110110", '1', '1', "11", "011", "110", "010", '0', '-', "00"), -- i=3328
      ("1011101000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3329
      ("0101001000110000", '0', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3330
      ("0101101000110000", '1', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3331
      ("0101101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3332
      ("0100001000110000", '0', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3333
      ("0100101000110000", '1', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3334
      ("0100101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3335
      ("0000001000010000", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3336
      ("0000101000010000", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3337
      ("0000101000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3338
      ("1000001000110111", '0', '1', "00", "011", "111", "010", '0', '-', "00"), -- i=3339
      ("1000101000110111", '1', '1', "00", "011", "111", "010", '0', '-', "00"), -- i=3340
      ("1000101000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3341
      ("1001001000110111", '0', '1', "01", "011", "111", "010", '0', '-', "00"), -- i=3342
      ("1001101000110111", '1', '1', "01", "011", "111", "010", '0', '-', "00"), -- i=3343
      ("1001101000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3344
      ("1010001000110111", '0', '1', "10", "011", "111", "010", '0', '-', "00"), -- i=3345
      ("1010101000110111", '1', '1', "10", "011", "111", "010", '0', '-', "00"), -- i=3346
      ("1010101000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3347
      ("1011001000110111", '0', '1', "11", "011", "111", "010", '0', '-', "00"), -- i=3348
      ("1011101000110111", '1', '1', "11", "011", "111", "010", '0', '-', "00"), -- i=3349
      ("1011101000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3350
      ("0101001000110000", '0', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3351
      ("0101101000110000", '1', '1', "--", "011", "---", "010", '0', '1', "01"), -- i=3352
      ("0101101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3353
      ("0100001000110000", '0', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3354
      ("0100101000110000", '1', '0', "--", "011", "010", "---", '1', '-', "--"), -- i=3355
      ("0100101000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3356
      ("0000001010000111", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3357
      ("0000101010000111", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3358
      ("0000101010000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3359
      ("1000001001000000", '0', '1', "00", "100", "000", "010", '0', '-', "00"), -- i=3360
      ("1000101001000000", '1', '1', "00", "100", "000", "010", '0', '-', "00"), -- i=3361
      ("1000101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3362
      ("1001001001000000", '0', '1', "01", "100", "000", "010", '0', '-', "00"), -- i=3363
      ("1001101001000000", '1', '1', "01", "100", "000", "010", '0', '-', "00"), -- i=3364
      ("1001101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3365
      ("1010001001000000", '0', '1', "10", "100", "000", "010", '0', '-', "00"), -- i=3366
      ("1010101001000000", '1', '1', "10", "100", "000", "010", '0', '-', "00"), -- i=3367
      ("1010101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3368
      ("1011001001000000", '0', '1', "11", "100", "000", "010", '0', '-', "00"), -- i=3369
      ("1011101001000000", '1', '1', "11", "100", "000", "010", '0', '-', "00"), -- i=3370
      ("1011101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3371
      ("0101001001000000", '0', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3372
      ("0101101001000000", '1', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3373
      ("0101101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3374
      ("0100001001000000", '0', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3375
      ("0100101001000000", '1', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3376
      ("0100101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3377
      ("0000001010101000", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3378
      ("0000101010101000", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3379
      ("0000101010101000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3380
      ("1000001001000001", '0', '1', "00", "100", "001", "010", '0', '-', "00"), -- i=3381
      ("1000101001000001", '1', '1', "00", "100", "001", "010", '0', '-', "00"), -- i=3382
      ("1000101001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3383
      ("1001001001000001", '0', '1', "01", "100", "001", "010", '0', '-', "00"), -- i=3384
      ("1001101001000001", '1', '1', "01", "100", "001", "010", '0', '-', "00"), -- i=3385
      ("1001101001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3386
      ("1010001001000001", '0', '1', "10", "100", "001", "010", '0', '-', "00"), -- i=3387
      ("1010101001000001", '1', '1', "10", "100", "001", "010", '0', '-', "00"), -- i=3388
      ("1010101001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3389
      ("1011001001000001", '0', '1', "11", "100", "001", "010", '0', '-', "00"), -- i=3390
      ("1011101001000001", '1', '1', "11", "100", "001", "010", '0', '-', "00"), -- i=3391
      ("1011101001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3392
      ("0101001001000000", '0', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3393
      ("0101101001000000", '1', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3394
      ("0101101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3395
      ("0100001001000000", '0', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3396
      ("0100101001000000", '1', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3397
      ("0100101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3398
      ("0000001010010101", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3399
      ("0000101010010101", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3400
      ("0000101010010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3401
      ("1000001001000010", '0', '1', "00", "100", "010", "010", '0', '-', "00"), -- i=3402
      ("1000101001000010", '1', '1', "00", "100", "010", "010", '0', '-', "00"), -- i=3403
      ("1000101001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3404
      ("1001001001000010", '0', '1', "01", "100", "010", "010", '0', '-', "00"), -- i=3405
      ("1001101001000010", '1', '1', "01", "100", "010", "010", '0', '-', "00"), -- i=3406
      ("1001101001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3407
      ("1010001001000010", '0', '1', "10", "100", "010", "010", '0', '-', "00"), -- i=3408
      ("1010101001000010", '1', '1', "10", "100", "010", "010", '0', '-', "00"), -- i=3409
      ("1010101001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3410
      ("1011001001000010", '0', '1', "11", "100", "010", "010", '0', '-', "00"), -- i=3411
      ("1011101001000010", '1', '1', "11", "100", "010", "010", '0', '-', "00"), -- i=3412
      ("1011101001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3413
      ("0101001001000000", '0', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3414
      ("0101101001000000", '1', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3415
      ("0101101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3416
      ("0100001001000000", '0', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3417
      ("0100101001000000", '1', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3418
      ("0100101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3419
      ("0000001000011111", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3420
      ("0000101000011111", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3421
      ("0000101000011111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3422
      ("1000001001000011", '0', '1', "00", "100", "011", "010", '0', '-', "00"), -- i=3423
      ("1000101001000011", '1', '1', "00", "100", "011", "010", '0', '-', "00"), -- i=3424
      ("1000101001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3425
      ("1001001001000011", '0', '1', "01", "100", "011", "010", '0', '-', "00"), -- i=3426
      ("1001101001000011", '1', '1', "01", "100", "011", "010", '0', '-', "00"), -- i=3427
      ("1001101001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3428
      ("1010001001000011", '0', '1', "10", "100", "011", "010", '0', '-', "00"), -- i=3429
      ("1010101001000011", '1', '1', "10", "100", "011", "010", '0', '-', "00"), -- i=3430
      ("1010101001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3431
      ("1011001001000011", '0', '1', "11", "100", "011", "010", '0', '-', "00"), -- i=3432
      ("1011101001000011", '1', '1', "11", "100", "011", "010", '0', '-', "00"), -- i=3433
      ("1011101001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3434
      ("0101001001000000", '0', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3435
      ("0101101001000000", '1', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3436
      ("0101101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3437
      ("0100001001000000", '0', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3438
      ("0100101001000000", '1', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3439
      ("0100101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3440
      ("0000001000010101", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3441
      ("0000101000010101", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3442
      ("0000101000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3443
      ("1000001001000100", '0', '1', "00", "100", "100", "010", '0', '-', "00"), -- i=3444
      ("1000101001000100", '1', '1', "00", "100", "100", "010", '0', '-', "00"), -- i=3445
      ("1000101001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3446
      ("1001001001000100", '0', '1', "01", "100", "100", "010", '0', '-', "00"), -- i=3447
      ("1001101001000100", '1', '1', "01", "100", "100", "010", '0', '-', "00"), -- i=3448
      ("1001101001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3449
      ("1010001001000100", '0', '1', "10", "100", "100", "010", '0', '-', "00"), -- i=3450
      ("1010101001000100", '1', '1', "10", "100", "100", "010", '0', '-', "00"), -- i=3451
      ("1010101001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3452
      ("1011001001000100", '0', '1', "11", "100", "100", "010", '0', '-', "00"), -- i=3453
      ("1011101001000100", '1', '1', "11", "100", "100", "010", '0', '-', "00"), -- i=3454
      ("1011101001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3455
      ("0101001001000000", '0', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3456
      ("0101101001000000", '1', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3457
      ("0101101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3458
      ("0100001001000000", '0', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3459
      ("0100101001000000", '1', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3460
      ("0100101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3461
      ("0000001001001000", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3462
      ("0000101001001000", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3463
      ("0000101001001000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3464
      ("1000001001000101", '0', '1', "00", "100", "101", "010", '0', '-', "00"), -- i=3465
      ("1000101001000101", '1', '1', "00", "100", "101", "010", '0', '-', "00"), -- i=3466
      ("1000101001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3467
      ("1001001001000101", '0', '1', "01", "100", "101", "010", '0', '-', "00"), -- i=3468
      ("1001101001000101", '1', '1', "01", "100", "101", "010", '0', '-', "00"), -- i=3469
      ("1001101001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3470
      ("1010001001000101", '0', '1', "10", "100", "101", "010", '0', '-', "00"), -- i=3471
      ("1010101001000101", '1', '1', "10", "100", "101", "010", '0', '-', "00"), -- i=3472
      ("1010101001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3473
      ("1011001001000101", '0', '1', "11", "100", "101", "010", '0', '-', "00"), -- i=3474
      ("1011101001000101", '1', '1', "11", "100", "101", "010", '0', '-', "00"), -- i=3475
      ("1011101001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3476
      ("0101001001000000", '0', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3477
      ("0101101001000000", '1', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3478
      ("0101101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3479
      ("0100001001000000", '0', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3480
      ("0100101001000000", '1', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3481
      ("0100101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3482
      ("0000001000111100", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3483
      ("0000101000111100", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3484
      ("0000101000111100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3485
      ("1000001001000110", '0', '1', "00", "100", "110", "010", '0', '-', "00"), -- i=3486
      ("1000101001000110", '1', '1', "00", "100", "110", "010", '0', '-', "00"), -- i=3487
      ("1000101001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3488
      ("1001001001000110", '0', '1', "01", "100", "110", "010", '0', '-', "00"), -- i=3489
      ("1001101001000110", '1', '1', "01", "100", "110", "010", '0', '-', "00"), -- i=3490
      ("1001101001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3491
      ("1010001001000110", '0', '1', "10", "100", "110", "010", '0', '-', "00"), -- i=3492
      ("1010101001000110", '1', '1', "10", "100", "110", "010", '0', '-', "00"), -- i=3493
      ("1010101001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3494
      ("1011001001000110", '0', '1', "11", "100", "110", "010", '0', '-', "00"), -- i=3495
      ("1011101001000110", '1', '1', "11", "100", "110", "010", '0', '-', "00"), -- i=3496
      ("1011101001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3497
      ("0101001001000000", '0', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3498
      ("0101101001000000", '1', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3499
      ("0101101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3500
      ("0100001001000000", '0', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3501
      ("0100101001000000", '1', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3502
      ("0100101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3503
      ("0000001011011010", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3504
      ("0000101011011010", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3505
      ("0000101011011010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3506
      ("1000001001000111", '0', '1', "00", "100", "111", "010", '0', '-', "00"), -- i=3507
      ("1000101001000111", '1', '1', "00", "100", "111", "010", '0', '-', "00"), -- i=3508
      ("1000101001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3509
      ("1001001001000111", '0', '1', "01", "100", "111", "010", '0', '-', "00"), -- i=3510
      ("1001101001000111", '1', '1', "01", "100", "111", "010", '0', '-', "00"), -- i=3511
      ("1001101001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3512
      ("1010001001000111", '0', '1', "10", "100", "111", "010", '0', '-', "00"), -- i=3513
      ("1010101001000111", '1', '1', "10", "100", "111", "010", '0', '-', "00"), -- i=3514
      ("1010101001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3515
      ("1011001001000111", '0', '1', "11", "100", "111", "010", '0', '-', "00"), -- i=3516
      ("1011101001000111", '1', '1', "11", "100", "111", "010", '0', '-', "00"), -- i=3517
      ("1011101001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3518
      ("0101001001000000", '0', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3519
      ("0101101001000000", '1', '1', "--", "100", "---", "010", '0', '1', "01"), -- i=3520
      ("0101101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3521
      ("0100001001000000", '0', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3522
      ("0100101001000000", '1', '0', "--", "100", "010", "---", '1', '-', "--"), -- i=3523
      ("0100101001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3524
      ("0000001001001000", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3525
      ("0000101001001000", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3526
      ("0000101001001000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3527
      ("1000001001010000", '0', '1', "00", "101", "000", "010", '0', '-', "00"), -- i=3528
      ("1000101001010000", '1', '1', "00", "101", "000", "010", '0', '-', "00"), -- i=3529
      ("1000101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3530
      ("1001001001010000", '0', '1', "01", "101", "000", "010", '0', '-', "00"), -- i=3531
      ("1001101001010000", '1', '1', "01", "101", "000", "010", '0', '-', "00"), -- i=3532
      ("1001101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3533
      ("1010001001010000", '0', '1', "10", "101", "000", "010", '0', '-', "00"), -- i=3534
      ("1010101001010000", '1', '1', "10", "101", "000", "010", '0', '-', "00"), -- i=3535
      ("1010101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3536
      ("1011001001010000", '0', '1', "11", "101", "000", "010", '0', '-', "00"), -- i=3537
      ("1011101001010000", '1', '1', "11", "101", "000", "010", '0', '-', "00"), -- i=3538
      ("1011101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3539
      ("0101001001010000", '0', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3540
      ("0101101001010000", '1', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3541
      ("0101101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3542
      ("0100001001010000", '0', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3543
      ("0100101001010000", '1', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3544
      ("0100101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3545
      ("0000001011101001", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3546
      ("0000101011101001", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3547
      ("0000101011101001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3548
      ("1000001001010001", '0', '1', "00", "101", "001", "010", '0', '-', "00"), -- i=3549
      ("1000101001010001", '1', '1', "00", "101", "001", "010", '0', '-', "00"), -- i=3550
      ("1000101001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3551
      ("1001001001010001", '0', '1', "01", "101", "001", "010", '0', '-', "00"), -- i=3552
      ("1001101001010001", '1', '1', "01", "101", "001", "010", '0', '-', "00"), -- i=3553
      ("1001101001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3554
      ("1010001001010001", '0', '1', "10", "101", "001", "010", '0', '-', "00"), -- i=3555
      ("1010101001010001", '1', '1', "10", "101", "001", "010", '0', '-', "00"), -- i=3556
      ("1010101001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3557
      ("1011001001010001", '0', '1', "11", "101", "001", "010", '0', '-', "00"), -- i=3558
      ("1011101001010001", '1', '1', "11", "101", "001", "010", '0', '-', "00"), -- i=3559
      ("1011101001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3560
      ("0101001001010000", '0', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3561
      ("0101101001010000", '1', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3562
      ("0101101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3563
      ("0100001001010000", '0', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3564
      ("0100101001010000", '1', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3565
      ("0100101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3566
      ("0000001010111000", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3567
      ("0000101010111000", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3568
      ("0000101010111000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3569
      ("1000001001010010", '0', '1', "00", "101", "010", "010", '0', '-', "00"), -- i=3570
      ("1000101001010010", '1', '1', "00", "101", "010", "010", '0', '-', "00"), -- i=3571
      ("1000101001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3572
      ("1001001001010010", '0', '1', "01", "101", "010", "010", '0', '-', "00"), -- i=3573
      ("1001101001010010", '1', '1', "01", "101", "010", "010", '0', '-', "00"), -- i=3574
      ("1001101001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3575
      ("1010001001010010", '0', '1', "10", "101", "010", "010", '0', '-', "00"), -- i=3576
      ("1010101001010010", '1', '1', "10", "101", "010", "010", '0', '-', "00"), -- i=3577
      ("1010101001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3578
      ("1011001001010010", '0', '1', "11", "101", "010", "010", '0', '-', "00"), -- i=3579
      ("1011101001010010", '1', '1', "11", "101", "010", "010", '0', '-', "00"), -- i=3580
      ("1011101001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3581
      ("0101001001010000", '0', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3582
      ("0101101001010000", '1', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3583
      ("0101101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3584
      ("0100001001010000", '0', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3585
      ("0100101001010000", '1', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3586
      ("0100101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3587
      ("0000001010000110", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3588
      ("0000101010000110", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3589
      ("0000101010000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3590
      ("1000001001010011", '0', '1', "00", "101", "011", "010", '0', '-', "00"), -- i=3591
      ("1000101001010011", '1', '1', "00", "101", "011", "010", '0', '-', "00"), -- i=3592
      ("1000101001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3593
      ("1001001001010011", '0', '1', "01", "101", "011", "010", '0', '-', "00"), -- i=3594
      ("1001101001010011", '1', '1', "01", "101", "011", "010", '0', '-', "00"), -- i=3595
      ("1001101001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3596
      ("1010001001010011", '0', '1', "10", "101", "011", "010", '0', '-', "00"), -- i=3597
      ("1010101001010011", '1', '1', "10", "101", "011", "010", '0', '-', "00"), -- i=3598
      ("1010101001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3599
      ("1011001001010011", '0', '1', "11", "101", "011", "010", '0', '-', "00"), -- i=3600
      ("1011101001010011", '1', '1', "11", "101", "011", "010", '0', '-', "00"), -- i=3601
      ("1011101001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3602
      ("0101001001010000", '0', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3603
      ("0101101001010000", '1', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3604
      ("0101101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3605
      ("0100001001010000", '0', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3606
      ("0100101001010000", '1', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3607
      ("0100101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3608
      ("0000001011110001", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3609
      ("0000101011110001", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3610
      ("0000101011110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3611
      ("1000001001010100", '0', '1', "00", "101", "100", "010", '0', '-', "00"), -- i=3612
      ("1000101001010100", '1', '1', "00", "101", "100", "010", '0', '-', "00"), -- i=3613
      ("1000101001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3614
      ("1001001001010100", '0', '1', "01", "101", "100", "010", '0', '-', "00"), -- i=3615
      ("1001101001010100", '1', '1', "01", "101", "100", "010", '0', '-', "00"), -- i=3616
      ("1001101001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3617
      ("1010001001010100", '0', '1', "10", "101", "100", "010", '0', '-', "00"), -- i=3618
      ("1010101001010100", '1', '1', "10", "101", "100", "010", '0', '-', "00"), -- i=3619
      ("1010101001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3620
      ("1011001001010100", '0', '1', "11", "101", "100", "010", '0', '-', "00"), -- i=3621
      ("1011101001010100", '1', '1', "11", "101", "100", "010", '0', '-', "00"), -- i=3622
      ("1011101001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3623
      ("0101001001010000", '0', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3624
      ("0101101001010000", '1', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3625
      ("0101101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3626
      ("0100001001010000", '0', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3627
      ("0100101001010000", '1', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3628
      ("0100101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3629
      ("0000001010100000", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3630
      ("0000101010100000", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3631
      ("0000101010100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3632
      ("1000001001010101", '0', '1', "00", "101", "101", "010", '0', '-', "00"), -- i=3633
      ("1000101001010101", '1', '1', "00", "101", "101", "010", '0', '-', "00"), -- i=3634
      ("1000101001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3635
      ("1001001001010101", '0', '1', "01", "101", "101", "010", '0', '-', "00"), -- i=3636
      ("1001101001010101", '1', '1', "01", "101", "101", "010", '0', '-', "00"), -- i=3637
      ("1001101001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3638
      ("1010001001010101", '0', '1', "10", "101", "101", "010", '0', '-', "00"), -- i=3639
      ("1010101001010101", '1', '1', "10", "101", "101", "010", '0', '-', "00"), -- i=3640
      ("1010101001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3641
      ("1011001001010101", '0', '1', "11", "101", "101", "010", '0', '-', "00"), -- i=3642
      ("1011101001010101", '1', '1', "11", "101", "101", "010", '0', '-', "00"), -- i=3643
      ("1011101001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3644
      ("0101001001010000", '0', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3645
      ("0101101001010000", '1', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3646
      ("0101101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3647
      ("0100001001010000", '0', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3648
      ("0100101001010000", '1', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3649
      ("0100101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3650
      ("0000001010110100", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3651
      ("0000101010110100", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3652
      ("0000101010110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3653
      ("1000001001010110", '0', '1', "00", "101", "110", "010", '0', '-', "00"), -- i=3654
      ("1000101001010110", '1', '1', "00", "101", "110", "010", '0', '-', "00"), -- i=3655
      ("1000101001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3656
      ("1001001001010110", '0', '1', "01", "101", "110", "010", '0', '-', "00"), -- i=3657
      ("1001101001010110", '1', '1', "01", "101", "110", "010", '0', '-', "00"), -- i=3658
      ("1001101001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3659
      ("1010001001010110", '0', '1', "10", "101", "110", "010", '0', '-', "00"), -- i=3660
      ("1010101001010110", '1', '1', "10", "101", "110", "010", '0', '-', "00"), -- i=3661
      ("1010101001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3662
      ("1011001001010110", '0', '1', "11", "101", "110", "010", '0', '-', "00"), -- i=3663
      ("1011101001010110", '1', '1', "11", "101", "110", "010", '0', '-', "00"), -- i=3664
      ("1011101001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3665
      ("0101001001010000", '0', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3666
      ("0101101001010000", '1', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3667
      ("0101101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3668
      ("0100001001010000", '0', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3669
      ("0100101001010000", '1', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3670
      ("0100101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3671
      ("0000001010000111", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3672
      ("0000101010000111", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3673
      ("0000101010000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3674
      ("1000001001010111", '0', '1', "00", "101", "111", "010", '0', '-', "00"), -- i=3675
      ("1000101001010111", '1', '1', "00", "101", "111", "010", '0', '-', "00"), -- i=3676
      ("1000101001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3677
      ("1001001001010111", '0', '1', "01", "101", "111", "010", '0', '-', "00"), -- i=3678
      ("1001101001010111", '1', '1', "01", "101", "111", "010", '0', '-', "00"), -- i=3679
      ("1001101001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3680
      ("1010001001010111", '0', '1', "10", "101", "111", "010", '0', '-', "00"), -- i=3681
      ("1010101001010111", '1', '1', "10", "101", "111", "010", '0', '-', "00"), -- i=3682
      ("1010101001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3683
      ("1011001001010111", '0', '1', "11", "101", "111", "010", '0', '-', "00"), -- i=3684
      ("1011101001010111", '1', '1', "11", "101", "111", "010", '0', '-', "00"), -- i=3685
      ("1011101001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3686
      ("0101001001010000", '0', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3687
      ("0101101001010000", '1', '1', "--", "101", "---", "010", '0', '1', "01"), -- i=3688
      ("0101101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3689
      ("0100001001010000", '0', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3690
      ("0100101001010000", '1', '0', "--", "101", "010", "---", '1', '-', "--"), -- i=3691
      ("0100101001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3692
      ("0000001010101011", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3693
      ("0000101010101011", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3694
      ("0000101010101011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3695
      ("1000001001100000", '0', '1', "00", "110", "000", "010", '0', '-', "00"), -- i=3696
      ("1000101001100000", '1', '1', "00", "110", "000", "010", '0', '-', "00"), -- i=3697
      ("1000101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3698
      ("1001001001100000", '0', '1', "01", "110", "000", "010", '0', '-', "00"), -- i=3699
      ("1001101001100000", '1', '1', "01", "110", "000", "010", '0', '-', "00"), -- i=3700
      ("1001101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3701
      ("1010001001100000", '0', '1', "10", "110", "000", "010", '0', '-', "00"), -- i=3702
      ("1010101001100000", '1', '1', "10", "110", "000", "010", '0', '-', "00"), -- i=3703
      ("1010101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3704
      ("1011001001100000", '0', '1', "11", "110", "000", "010", '0', '-', "00"), -- i=3705
      ("1011101001100000", '1', '1', "11", "110", "000", "010", '0', '-', "00"), -- i=3706
      ("1011101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3707
      ("0101001001100000", '0', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3708
      ("0101101001100000", '1', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3709
      ("0101101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3710
      ("0100001001100000", '0', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3711
      ("0100101001100000", '1', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3712
      ("0100101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3713
      ("0000001011010110", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3714
      ("0000101011010110", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3715
      ("0000101011010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3716
      ("1000001001100001", '0', '1', "00", "110", "001", "010", '0', '-', "00"), -- i=3717
      ("1000101001100001", '1', '1', "00", "110", "001", "010", '0', '-', "00"), -- i=3718
      ("1000101001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3719
      ("1001001001100001", '0', '1', "01", "110", "001", "010", '0', '-', "00"), -- i=3720
      ("1001101001100001", '1', '1', "01", "110", "001", "010", '0', '-', "00"), -- i=3721
      ("1001101001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3722
      ("1010001001100001", '0', '1', "10", "110", "001", "010", '0', '-', "00"), -- i=3723
      ("1010101001100001", '1', '1', "10", "110", "001", "010", '0', '-', "00"), -- i=3724
      ("1010101001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3725
      ("1011001001100001", '0', '1', "11", "110", "001", "010", '0', '-', "00"), -- i=3726
      ("1011101001100001", '1', '1', "11", "110", "001", "010", '0', '-', "00"), -- i=3727
      ("1011101001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3728
      ("0101001001100000", '0', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3729
      ("0101101001100000", '1', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3730
      ("0101101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3731
      ("0100001001100000", '0', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3732
      ("0100101001100000", '1', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3733
      ("0100101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3734
      ("0000001000001100", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3735
      ("0000101000001100", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3736
      ("0000101000001100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3737
      ("1000001001100010", '0', '1', "00", "110", "010", "010", '0', '-', "00"), -- i=3738
      ("1000101001100010", '1', '1', "00", "110", "010", "010", '0', '-', "00"), -- i=3739
      ("1000101001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3740
      ("1001001001100010", '0', '1', "01", "110", "010", "010", '0', '-', "00"), -- i=3741
      ("1001101001100010", '1', '1', "01", "110", "010", "010", '0', '-', "00"), -- i=3742
      ("1001101001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3743
      ("1010001001100010", '0', '1', "10", "110", "010", "010", '0', '-', "00"), -- i=3744
      ("1010101001100010", '1', '1', "10", "110", "010", "010", '0', '-', "00"), -- i=3745
      ("1010101001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3746
      ("1011001001100010", '0', '1', "11", "110", "010", "010", '0', '-', "00"), -- i=3747
      ("1011101001100010", '1', '1', "11", "110", "010", "010", '0', '-', "00"), -- i=3748
      ("1011101001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3749
      ("0101001001100000", '0', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3750
      ("0101101001100000", '1', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3751
      ("0101101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3752
      ("0100001001100000", '0', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3753
      ("0100101001100000", '1', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3754
      ("0100101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3755
      ("0000001010111100", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3756
      ("0000101010111100", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3757
      ("0000101010111100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3758
      ("1000001001100011", '0', '1', "00", "110", "011", "010", '0', '-', "00"), -- i=3759
      ("1000101001100011", '1', '1', "00", "110", "011", "010", '0', '-', "00"), -- i=3760
      ("1000101001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3761
      ("1001001001100011", '0', '1', "01", "110", "011", "010", '0', '-', "00"), -- i=3762
      ("1001101001100011", '1', '1', "01", "110", "011", "010", '0', '-', "00"), -- i=3763
      ("1001101001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3764
      ("1010001001100011", '0', '1', "10", "110", "011", "010", '0', '-', "00"), -- i=3765
      ("1010101001100011", '1', '1', "10", "110", "011", "010", '0', '-', "00"), -- i=3766
      ("1010101001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3767
      ("1011001001100011", '0', '1', "11", "110", "011", "010", '0', '-', "00"), -- i=3768
      ("1011101001100011", '1', '1', "11", "110", "011", "010", '0', '-', "00"), -- i=3769
      ("1011101001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3770
      ("0101001001100000", '0', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3771
      ("0101101001100000", '1', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3772
      ("0101101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3773
      ("0100001001100000", '0', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3774
      ("0100101001100000", '1', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3775
      ("0100101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3776
      ("0000001001010011", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3777
      ("0000101001010011", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3778
      ("0000101001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3779
      ("1000001001100100", '0', '1', "00", "110", "100", "010", '0', '-', "00"), -- i=3780
      ("1000101001100100", '1', '1', "00", "110", "100", "010", '0', '-', "00"), -- i=3781
      ("1000101001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3782
      ("1001001001100100", '0', '1', "01", "110", "100", "010", '0', '-', "00"), -- i=3783
      ("1001101001100100", '1', '1', "01", "110", "100", "010", '0', '-', "00"), -- i=3784
      ("1001101001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3785
      ("1010001001100100", '0', '1', "10", "110", "100", "010", '0', '-', "00"), -- i=3786
      ("1010101001100100", '1', '1', "10", "110", "100", "010", '0', '-', "00"), -- i=3787
      ("1010101001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3788
      ("1011001001100100", '0', '1', "11", "110", "100", "010", '0', '-', "00"), -- i=3789
      ("1011101001100100", '1', '1', "11", "110", "100", "010", '0', '-', "00"), -- i=3790
      ("1011101001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3791
      ("0101001001100000", '0', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3792
      ("0101101001100000", '1', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3793
      ("0101101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3794
      ("0100001001100000", '0', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3795
      ("0100101001100000", '1', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3796
      ("0100101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3797
      ("0000001001000111", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3798
      ("0000101001000111", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3799
      ("0000101001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3800
      ("1000001001100101", '0', '1', "00", "110", "101", "010", '0', '-', "00"), -- i=3801
      ("1000101001100101", '1', '1', "00", "110", "101", "010", '0', '-', "00"), -- i=3802
      ("1000101001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3803
      ("1001001001100101", '0', '1', "01", "110", "101", "010", '0', '-', "00"), -- i=3804
      ("1001101001100101", '1', '1', "01", "110", "101", "010", '0', '-', "00"), -- i=3805
      ("1001101001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3806
      ("1010001001100101", '0', '1', "10", "110", "101", "010", '0', '-', "00"), -- i=3807
      ("1010101001100101", '1', '1', "10", "110", "101", "010", '0', '-', "00"), -- i=3808
      ("1010101001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3809
      ("1011001001100101", '0', '1', "11", "110", "101", "010", '0', '-', "00"), -- i=3810
      ("1011101001100101", '1', '1', "11", "110", "101", "010", '0', '-', "00"), -- i=3811
      ("1011101001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3812
      ("0101001001100000", '0', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3813
      ("0101101001100000", '1', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3814
      ("0101101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3815
      ("0100001001100000", '0', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3816
      ("0100101001100000", '1', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3817
      ("0100101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3818
      ("0000001011011011", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3819
      ("0000101011011011", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3820
      ("0000101011011011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3821
      ("1000001001100110", '0', '1', "00", "110", "110", "010", '0', '-', "00"), -- i=3822
      ("1000101001100110", '1', '1', "00", "110", "110", "010", '0', '-', "00"), -- i=3823
      ("1000101001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3824
      ("1001001001100110", '0', '1', "01", "110", "110", "010", '0', '-', "00"), -- i=3825
      ("1001101001100110", '1', '1', "01", "110", "110", "010", '0', '-', "00"), -- i=3826
      ("1001101001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3827
      ("1010001001100110", '0', '1', "10", "110", "110", "010", '0', '-', "00"), -- i=3828
      ("1010101001100110", '1', '1', "10", "110", "110", "010", '0', '-', "00"), -- i=3829
      ("1010101001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3830
      ("1011001001100110", '0', '1', "11", "110", "110", "010", '0', '-', "00"), -- i=3831
      ("1011101001100110", '1', '1', "11", "110", "110", "010", '0', '-', "00"), -- i=3832
      ("1011101001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3833
      ("0101001001100000", '0', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3834
      ("0101101001100000", '1', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3835
      ("0101101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3836
      ("0100001001100000", '0', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3837
      ("0100101001100000", '1', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3838
      ("0100101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3839
      ("0000001000101100", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3840
      ("0000101000101100", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3841
      ("0000101000101100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3842
      ("1000001001100111", '0', '1', "00", "110", "111", "010", '0', '-', "00"), -- i=3843
      ("1000101001100111", '1', '1', "00", "110", "111", "010", '0', '-', "00"), -- i=3844
      ("1000101001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3845
      ("1001001001100111", '0', '1', "01", "110", "111", "010", '0', '-', "00"), -- i=3846
      ("1001101001100111", '1', '1', "01", "110", "111", "010", '0', '-', "00"), -- i=3847
      ("1001101001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3848
      ("1010001001100111", '0', '1', "10", "110", "111", "010", '0', '-', "00"), -- i=3849
      ("1010101001100111", '1', '1', "10", "110", "111", "010", '0', '-', "00"), -- i=3850
      ("1010101001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3851
      ("1011001001100111", '0', '1', "11", "110", "111", "010", '0', '-', "00"), -- i=3852
      ("1011101001100111", '1', '1', "11", "110", "111", "010", '0', '-', "00"), -- i=3853
      ("1011101001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3854
      ("0101001001100000", '0', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3855
      ("0101101001100000", '1', '1', "--", "110", "---", "010", '0', '1', "01"), -- i=3856
      ("0101101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3857
      ("0100001001100000", '0', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3858
      ("0100101001100000", '1', '0', "--", "110", "010", "---", '1', '-', "--"), -- i=3859
      ("0100101001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3860
      ("0000001011111011", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3861
      ("0000101011111011", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3862
      ("0000101011111011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3863
      ("1000001001110000", '0', '1', "00", "111", "000", "010", '0', '-', "00"), -- i=3864
      ("1000101001110000", '1', '1', "00", "111", "000", "010", '0', '-', "00"), -- i=3865
      ("1000101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3866
      ("1001001001110000", '0', '1', "01", "111", "000", "010", '0', '-', "00"), -- i=3867
      ("1001101001110000", '1', '1', "01", "111", "000", "010", '0', '-', "00"), -- i=3868
      ("1001101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3869
      ("1010001001110000", '0', '1', "10", "111", "000", "010", '0', '-', "00"), -- i=3870
      ("1010101001110000", '1', '1', "10", "111", "000", "010", '0', '-', "00"), -- i=3871
      ("1010101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3872
      ("1011001001110000", '0', '1', "11", "111", "000", "010", '0', '-', "00"), -- i=3873
      ("1011101001110000", '1', '1', "11", "111", "000", "010", '0', '-', "00"), -- i=3874
      ("1011101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3875
      ("0101001001110000", '0', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=3876
      ("0101101001110000", '1', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=3877
      ("0101101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3878
      ("0100001001110000", '0', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=3879
      ("0100101001110000", '1', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=3880
      ("0100101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3881
      ("0000001001000111", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3882
      ("0000101001000111", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3883
      ("0000101001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3884
      ("1000001001110001", '0', '1', "00", "111", "001", "010", '0', '-', "00"), -- i=3885
      ("1000101001110001", '1', '1', "00", "111", "001", "010", '0', '-', "00"), -- i=3886
      ("1000101001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3887
      ("1001001001110001", '0', '1', "01", "111", "001", "010", '0', '-', "00"), -- i=3888
      ("1001101001110001", '1', '1', "01", "111", "001", "010", '0', '-', "00"), -- i=3889
      ("1001101001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3890
      ("1010001001110001", '0', '1', "10", "111", "001", "010", '0', '-', "00"), -- i=3891
      ("1010101001110001", '1', '1', "10", "111", "001", "010", '0', '-', "00"), -- i=3892
      ("1010101001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3893
      ("1011001001110001", '0', '1', "11", "111", "001", "010", '0', '-', "00"), -- i=3894
      ("1011101001110001", '1', '1', "11", "111", "001", "010", '0', '-', "00"), -- i=3895
      ("1011101001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3896
      ("0101001001110000", '0', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=3897
      ("0101101001110000", '1', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=3898
      ("0101101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3899
      ("0100001001110000", '0', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=3900
      ("0100101001110000", '1', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=3901
      ("0100101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3902
      ("0000001000110100", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3903
      ("0000101000110100", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3904
      ("0000101000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3905
      ("1000001001110010", '0', '1', "00", "111", "010", "010", '0', '-', "00"), -- i=3906
      ("1000101001110010", '1', '1', "00", "111", "010", "010", '0', '-', "00"), -- i=3907
      ("1000101001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3908
      ("1001001001110010", '0', '1', "01", "111", "010", "010", '0', '-', "00"), -- i=3909
      ("1001101001110010", '1', '1', "01", "111", "010", "010", '0', '-', "00"), -- i=3910
      ("1001101001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3911
      ("1010001001110010", '0', '1', "10", "111", "010", "010", '0', '-', "00"), -- i=3912
      ("1010101001110010", '1', '1', "10", "111", "010", "010", '0', '-', "00"), -- i=3913
      ("1010101001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3914
      ("1011001001110010", '0', '1', "11", "111", "010", "010", '0', '-', "00"), -- i=3915
      ("1011101001110010", '1', '1', "11", "111", "010", "010", '0', '-', "00"), -- i=3916
      ("1011101001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3917
      ("0101001001110000", '0', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=3918
      ("0101101001110000", '1', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=3919
      ("0101101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3920
      ("0100001001110000", '0', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=3921
      ("0100101001110000", '1', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=3922
      ("0100101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3923
      ("0000001000111111", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3924
      ("0000101000111111", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3925
      ("0000101000111111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3926
      ("1000001001110011", '0', '1', "00", "111", "011", "010", '0', '-', "00"), -- i=3927
      ("1000101001110011", '1', '1', "00", "111", "011", "010", '0', '-', "00"), -- i=3928
      ("1000101001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3929
      ("1001001001110011", '0', '1', "01", "111", "011", "010", '0', '-', "00"), -- i=3930
      ("1001101001110011", '1', '1', "01", "111", "011", "010", '0', '-', "00"), -- i=3931
      ("1001101001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3932
      ("1010001001110011", '0', '1', "10", "111", "011", "010", '0', '-', "00"), -- i=3933
      ("1010101001110011", '1', '1', "10", "111", "011", "010", '0', '-', "00"), -- i=3934
      ("1010101001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3935
      ("1011001001110011", '0', '1', "11", "111", "011", "010", '0', '-', "00"), -- i=3936
      ("1011101001110011", '1', '1', "11", "111", "011", "010", '0', '-', "00"), -- i=3937
      ("1011101001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3938
      ("0101001001110000", '0', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=3939
      ("0101101001110000", '1', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=3940
      ("0101101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3941
      ("0100001001110000", '0', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=3942
      ("0100101001110000", '1', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=3943
      ("0100101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3944
      ("0000001001110111", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3945
      ("0000101001110111", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3946
      ("0000101001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3947
      ("1000001001110100", '0', '1', "00", "111", "100", "010", '0', '-', "00"), -- i=3948
      ("1000101001110100", '1', '1', "00", "111", "100", "010", '0', '-', "00"), -- i=3949
      ("1000101001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3950
      ("1001001001110100", '0', '1', "01", "111", "100", "010", '0', '-', "00"), -- i=3951
      ("1001101001110100", '1', '1', "01", "111", "100", "010", '0', '-', "00"), -- i=3952
      ("1001101001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3953
      ("1010001001110100", '0', '1', "10", "111", "100", "010", '0', '-', "00"), -- i=3954
      ("1010101001110100", '1', '1', "10", "111", "100", "010", '0', '-', "00"), -- i=3955
      ("1010101001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3956
      ("1011001001110100", '0', '1', "11", "111", "100", "010", '0', '-', "00"), -- i=3957
      ("1011101001110100", '1', '1', "11", "111", "100", "010", '0', '-', "00"), -- i=3958
      ("1011101001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3959
      ("0101001001110000", '0', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=3960
      ("0101101001110000", '1', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=3961
      ("0101101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3962
      ("0100001001110000", '0', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=3963
      ("0100101001110000", '1', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=3964
      ("0100101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3965
      ("0000001010000101", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3966
      ("0000101010000101", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3967
      ("0000101010000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3968
      ("1000001001110101", '0', '1', "00", "111", "101", "010", '0', '-', "00"), -- i=3969
      ("1000101001110101", '1', '1', "00", "111", "101", "010", '0', '-', "00"), -- i=3970
      ("1000101001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3971
      ("1001001001110101", '0', '1', "01", "111", "101", "010", '0', '-', "00"), -- i=3972
      ("1001101001110101", '1', '1', "01", "111", "101", "010", '0', '-', "00"), -- i=3973
      ("1001101001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3974
      ("1010001001110101", '0', '1', "10", "111", "101", "010", '0', '-', "00"), -- i=3975
      ("1010101001110101", '1', '1', "10", "111", "101", "010", '0', '-', "00"), -- i=3976
      ("1010101001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3977
      ("1011001001110101", '0', '1', "11", "111", "101", "010", '0', '-', "00"), -- i=3978
      ("1011101001110101", '1', '1', "11", "111", "101", "010", '0', '-', "00"), -- i=3979
      ("1011101001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3980
      ("0101001001110000", '0', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=3981
      ("0101101001110000", '1', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=3982
      ("0101101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3983
      ("0100001001110000", '0', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=3984
      ("0100101001110000", '1', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=3985
      ("0100101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3986
      ("0000001011100011", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3987
      ("0000101011100011", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=3988
      ("0000101011100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3989
      ("1000001001110110", '0', '1', "00", "111", "110", "010", '0', '-', "00"), -- i=3990
      ("1000101001110110", '1', '1', "00", "111", "110", "010", '0', '-', "00"), -- i=3991
      ("1000101001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3992
      ("1001001001110110", '0', '1', "01", "111", "110", "010", '0', '-', "00"), -- i=3993
      ("1001101001110110", '1', '1', "01", "111", "110", "010", '0', '-', "00"), -- i=3994
      ("1001101001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3995
      ("1010001001110110", '0', '1', "10", "111", "110", "010", '0', '-', "00"), -- i=3996
      ("1010101001110110", '1', '1', "10", "111", "110", "010", '0', '-', "00"), -- i=3997
      ("1010101001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=3998
      ("1011001001110110", '0', '1', "11", "111", "110", "010", '0', '-', "00"), -- i=3999
      ("1011101001110110", '1', '1', "11", "111", "110", "010", '0', '-', "00"), -- i=4000
      ("1011101001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4001
      ("0101001001110000", '0', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=4002
      ("0101101001110000", '1', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=4003
      ("0101101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4004
      ("0100001001110000", '0', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=4005
      ("0100101001110000", '1', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=4006
      ("0100101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4007
      ("0000001001101000", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=4008
      ("0000101001101000", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=4009
      ("0000101001101000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4010
      ("1000001001110111", '0', '1', "00", "111", "111", "010", '0', '-', "00"), -- i=4011
      ("1000101001110111", '1', '1', "00", "111", "111", "010", '0', '-', "00"), -- i=4012
      ("1000101001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4013
      ("1001001001110111", '0', '1', "01", "111", "111", "010", '0', '-', "00"), -- i=4014
      ("1001101001110111", '1', '1', "01", "111", "111", "010", '0', '-', "00"), -- i=4015
      ("1001101001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4016
      ("1010001001110111", '0', '1', "10", "111", "111", "010", '0', '-', "00"), -- i=4017
      ("1010101001110111", '1', '1', "10", "111", "111", "010", '0', '-', "00"), -- i=4018
      ("1010101001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4019
      ("1011001001110111", '0', '1', "11", "111", "111", "010", '0', '-', "00"), -- i=4020
      ("1011101001110111", '1', '1', "11", "111", "111", "010", '0', '-', "00"), -- i=4021
      ("1011101001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4022
      ("0101001001110000", '0', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=4023
      ("0101101001110000", '1', '1', "--", "111", "---", "010", '0', '1', "01"), -- i=4024
      ("0101101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4025
      ("0100001001110000", '0', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=4026
      ("0100101001110000", '1', '0', "--", "111", "010", "---", '1', '-', "--"), -- i=4027
      ("0100101001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4028
      ("0000001001000011", '0', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=4029
      ("0000101001000011", '1', '1', "--", "---", "---", "010", '0', '-', "10"), -- i=4030
      ("0000101001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4031
      ("1000001100000000", '0', '1', "00", "000", "000", "011", '0', '-', "00"), -- i=4032
      ("1000101100000000", '1', '1', "00", "000", "000", "011", '0', '-', "00"), -- i=4033
      ("1000101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4034
      ("1001001100000000", '0', '1', "01", "000", "000", "011", '0', '-', "00"), -- i=4035
      ("1001101100000000", '1', '1', "01", "000", "000", "011", '0', '-', "00"), -- i=4036
      ("1001101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4037
      ("1010001100000000", '0', '1', "10", "000", "000", "011", '0', '-', "00"), -- i=4038
      ("1010101100000000", '1', '1', "10", "000", "000", "011", '0', '-', "00"), -- i=4039
      ("1010101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4040
      ("1011001100000000", '0', '1', "11", "000", "000", "011", '0', '-', "00"), -- i=4041
      ("1011101100000000", '1', '1', "11", "000", "000", "011", '0', '-', "00"), -- i=4042
      ("1011101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4043
      ("0101001100000000", '0', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4044
      ("0101101100000000", '1', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4045
      ("0101101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4046
      ("0100001100000000", '0', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4047
      ("0100101100000000", '1', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4048
      ("0100101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4049
      ("0000001111000010", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4050
      ("0000101111000010", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4051
      ("0000101111000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4052
      ("1000001100000001", '0', '1', "00", "000", "001", "011", '0', '-', "00"), -- i=4053
      ("1000101100000001", '1', '1', "00", "000", "001", "011", '0', '-', "00"), -- i=4054
      ("1000101100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4055
      ("1001001100000001", '0', '1', "01", "000", "001", "011", '0', '-', "00"), -- i=4056
      ("1001101100000001", '1', '1', "01", "000", "001", "011", '0', '-', "00"), -- i=4057
      ("1001101100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4058
      ("1010001100000001", '0', '1', "10", "000", "001", "011", '0', '-', "00"), -- i=4059
      ("1010101100000001", '1', '1', "10", "000", "001", "011", '0', '-', "00"), -- i=4060
      ("1010101100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4061
      ("1011001100000001", '0', '1', "11", "000", "001", "011", '0', '-', "00"), -- i=4062
      ("1011101100000001", '1', '1', "11", "000", "001", "011", '0', '-', "00"), -- i=4063
      ("1011101100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4064
      ("0101001100000000", '0', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4065
      ("0101101100000000", '1', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4066
      ("0101101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4067
      ("0100001100000000", '0', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4068
      ("0100101100000000", '1', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4069
      ("0100101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4070
      ("0000001111000000", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4071
      ("0000101111000000", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4072
      ("0000101111000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4073
      ("1000001100000010", '0', '1', "00", "000", "010", "011", '0', '-', "00"), -- i=4074
      ("1000101100000010", '1', '1', "00", "000", "010", "011", '0', '-', "00"), -- i=4075
      ("1000101100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4076
      ("1001001100000010", '0', '1', "01", "000", "010", "011", '0', '-', "00"), -- i=4077
      ("1001101100000010", '1', '1', "01", "000", "010", "011", '0', '-', "00"), -- i=4078
      ("1001101100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4079
      ("1010001100000010", '0', '1', "10", "000", "010", "011", '0', '-', "00"), -- i=4080
      ("1010101100000010", '1', '1', "10", "000", "010", "011", '0', '-', "00"), -- i=4081
      ("1010101100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4082
      ("1011001100000010", '0', '1', "11", "000", "010", "011", '0', '-', "00"), -- i=4083
      ("1011101100000010", '1', '1', "11", "000", "010", "011", '0', '-', "00"), -- i=4084
      ("1011101100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4085
      ("0101001100000000", '0', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4086
      ("0101101100000000", '1', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4087
      ("0101101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4088
      ("0100001100000000", '0', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4089
      ("0100101100000000", '1', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4090
      ("0100101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4091
      ("0000001110010101", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4092
      ("0000101110010101", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4093
      ("0000101110010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4094
      ("1000001100000011", '0', '1', "00", "000", "011", "011", '0', '-', "00"), -- i=4095
      ("1000101100000011", '1', '1', "00", "000", "011", "011", '0', '-', "00"), -- i=4096
      ("1000101100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4097
      ("1001001100000011", '0', '1', "01", "000", "011", "011", '0', '-', "00"), -- i=4098
      ("1001101100000011", '1', '1', "01", "000", "011", "011", '0', '-', "00"), -- i=4099
      ("1001101100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4100
      ("1010001100000011", '0', '1', "10", "000", "011", "011", '0', '-', "00"), -- i=4101
      ("1010101100000011", '1', '1', "10", "000", "011", "011", '0', '-', "00"), -- i=4102
      ("1010101100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4103
      ("1011001100000011", '0', '1', "11", "000", "011", "011", '0', '-', "00"), -- i=4104
      ("1011101100000011", '1', '1', "11", "000", "011", "011", '0', '-', "00"), -- i=4105
      ("1011101100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4106
      ("0101001100000000", '0', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4107
      ("0101101100000000", '1', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4108
      ("0101101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4109
      ("0100001100000000", '0', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4110
      ("0100101100000000", '1', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4111
      ("0100101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4112
      ("0000001110001100", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4113
      ("0000101110001100", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4114
      ("0000101110001100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4115
      ("1000001100000100", '0', '1', "00", "000", "100", "011", '0', '-', "00"), -- i=4116
      ("1000101100000100", '1', '1', "00", "000", "100", "011", '0', '-', "00"), -- i=4117
      ("1000101100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4118
      ("1001001100000100", '0', '1', "01", "000", "100", "011", '0', '-', "00"), -- i=4119
      ("1001101100000100", '1', '1', "01", "000", "100", "011", '0', '-', "00"), -- i=4120
      ("1001101100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4121
      ("1010001100000100", '0', '1', "10", "000", "100", "011", '0', '-', "00"), -- i=4122
      ("1010101100000100", '1', '1', "10", "000", "100", "011", '0', '-', "00"), -- i=4123
      ("1010101100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4124
      ("1011001100000100", '0', '1', "11", "000", "100", "011", '0', '-', "00"), -- i=4125
      ("1011101100000100", '1', '1', "11", "000", "100", "011", '0', '-', "00"), -- i=4126
      ("1011101100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4127
      ("0101001100000000", '0', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4128
      ("0101101100000000", '1', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4129
      ("0101101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4130
      ("0100001100000000", '0', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4131
      ("0100101100000000", '1', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4132
      ("0100101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4133
      ("0000001111111000", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4134
      ("0000101111111000", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4135
      ("0000101111111000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4136
      ("1000001100000101", '0', '1', "00", "000", "101", "011", '0', '-', "00"), -- i=4137
      ("1000101100000101", '1', '1', "00", "000", "101", "011", '0', '-', "00"), -- i=4138
      ("1000101100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4139
      ("1001001100000101", '0', '1', "01", "000", "101", "011", '0', '-', "00"), -- i=4140
      ("1001101100000101", '1', '1', "01", "000", "101", "011", '0', '-', "00"), -- i=4141
      ("1001101100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4142
      ("1010001100000101", '0', '1', "10", "000", "101", "011", '0', '-', "00"), -- i=4143
      ("1010101100000101", '1', '1', "10", "000", "101", "011", '0', '-', "00"), -- i=4144
      ("1010101100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4145
      ("1011001100000101", '0', '1', "11", "000", "101", "011", '0', '-', "00"), -- i=4146
      ("1011101100000101", '1', '1', "11", "000", "101", "011", '0', '-', "00"), -- i=4147
      ("1011101100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4148
      ("0101001100000000", '0', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4149
      ("0101101100000000", '1', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4150
      ("0101101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4151
      ("0100001100000000", '0', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4152
      ("0100101100000000", '1', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4153
      ("0100101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4154
      ("0000001111101101", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4155
      ("0000101111101101", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4156
      ("0000101111101101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4157
      ("1000001100000110", '0', '1', "00", "000", "110", "011", '0', '-', "00"), -- i=4158
      ("1000101100000110", '1', '1', "00", "000", "110", "011", '0', '-', "00"), -- i=4159
      ("1000101100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4160
      ("1001001100000110", '0', '1', "01", "000", "110", "011", '0', '-', "00"), -- i=4161
      ("1001101100000110", '1', '1', "01", "000", "110", "011", '0', '-', "00"), -- i=4162
      ("1001101100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4163
      ("1010001100000110", '0', '1', "10", "000", "110", "011", '0', '-', "00"), -- i=4164
      ("1010101100000110", '1', '1', "10", "000", "110", "011", '0', '-', "00"), -- i=4165
      ("1010101100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4166
      ("1011001100000110", '0', '1', "11", "000", "110", "011", '0', '-', "00"), -- i=4167
      ("1011101100000110", '1', '1', "11", "000", "110", "011", '0', '-', "00"), -- i=4168
      ("1011101100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4169
      ("0101001100000000", '0', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4170
      ("0101101100000000", '1', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4171
      ("0101101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4172
      ("0100001100000000", '0', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4173
      ("0100101100000000", '1', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4174
      ("0100101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4175
      ("0000001100001110", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4176
      ("0000101100001110", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4177
      ("0000101100001110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4178
      ("1000001100000111", '0', '1', "00", "000", "111", "011", '0', '-', "00"), -- i=4179
      ("1000101100000111", '1', '1', "00", "000", "111", "011", '0', '-', "00"), -- i=4180
      ("1000101100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4181
      ("1001001100000111", '0', '1', "01", "000", "111", "011", '0', '-', "00"), -- i=4182
      ("1001101100000111", '1', '1', "01", "000", "111", "011", '0', '-', "00"), -- i=4183
      ("1001101100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4184
      ("1010001100000111", '0', '1', "10", "000", "111", "011", '0', '-', "00"), -- i=4185
      ("1010101100000111", '1', '1', "10", "000", "111", "011", '0', '-', "00"), -- i=4186
      ("1010101100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4187
      ("1011001100000111", '0', '1', "11", "000", "111", "011", '0', '-', "00"), -- i=4188
      ("1011101100000111", '1', '1', "11", "000", "111", "011", '0', '-', "00"), -- i=4189
      ("1011101100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4190
      ("0101001100000000", '0', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4191
      ("0101101100000000", '1', '1', "--", "000", "---", "011", '0', '1', "01"), -- i=4192
      ("0101101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4193
      ("0100001100000000", '0', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4194
      ("0100101100000000", '1', '0', "--", "000", "011", "---", '1', '-', "--"), -- i=4195
      ("0100101100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4196
      ("0000001111000111", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4197
      ("0000101111000111", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4198
      ("0000101111000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4199
      ("1000001100010000", '0', '1', "00", "001", "000", "011", '0', '-', "00"), -- i=4200
      ("1000101100010000", '1', '1', "00", "001", "000", "011", '0', '-', "00"), -- i=4201
      ("1000101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4202
      ("1001001100010000", '0', '1', "01", "001", "000", "011", '0', '-', "00"), -- i=4203
      ("1001101100010000", '1', '1', "01", "001", "000", "011", '0', '-', "00"), -- i=4204
      ("1001101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4205
      ("1010001100010000", '0', '1', "10", "001", "000", "011", '0', '-', "00"), -- i=4206
      ("1010101100010000", '1', '1', "10", "001", "000", "011", '0', '-', "00"), -- i=4207
      ("1010101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4208
      ("1011001100010000", '0', '1', "11", "001", "000", "011", '0', '-', "00"), -- i=4209
      ("1011101100010000", '1', '1', "11", "001", "000", "011", '0', '-', "00"), -- i=4210
      ("1011101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4211
      ("0101001100010000", '0', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4212
      ("0101101100010000", '1', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4213
      ("0101101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4214
      ("0100001100010000", '0', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4215
      ("0100101100010000", '1', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4216
      ("0100101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4217
      ("0000001100100110", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4218
      ("0000101100100110", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4219
      ("0000101100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4220
      ("1000001100010001", '0', '1', "00", "001", "001", "011", '0', '-', "00"), -- i=4221
      ("1000101100010001", '1', '1', "00", "001", "001", "011", '0', '-', "00"), -- i=4222
      ("1000101100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4223
      ("1001001100010001", '0', '1', "01", "001", "001", "011", '0', '-', "00"), -- i=4224
      ("1001101100010001", '1', '1', "01", "001", "001", "011", '0', '-', "00"), -- i=4225
      ("1001101100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4226
      ("1010001100010001", '0', '1', "10", "001", "001", "011", '0', '-', "00"), -- i=4227
      ("1010101100010001", '1', '1', "10", "001", "001", "011", '0', '-', "00"), -- i=4228
      ("1010101100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4229
      ("1011001100010001", '0', '1', "11", "001", "001", "011", '0', '-', "00"), -- i=4230
      ("1011101100010001", '1', '1', "11", "001", "001", "011", '0', '-', "00"), -- i=4231
      ("1011101100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4232
      ("0101001100010000", '0', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4233
      ("0101101100010000", '1', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4234
      ("0101101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4235
      ("0100001100010000", '0', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4236
      ("0100101100010000", '1', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4237
      ("0100101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4238
      ("0000001101110111", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4239
      ("0000101101110111", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4240
      ("0000101101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4241
      ("1000001100010010", '0', '1', "00", "001", "010", "011", '0', '-', "00"), -- i=4242
      ("1000101100010010", '1', '1', "00", "001", "010", "011", '0', '-', "00"), -- i=4243
      ("1000101100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4244
      ("1001001100010010", '0', '1', "01", "001", "010", "011", '0', '-', "00"), -- i=4245
      ("1001101100010010", '1', '1', "01", "001", "010", "011", '0', '-', "00"), -- i=4246
      ("1001101100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4247
      ("1010001100010010", '0', '1', "10", "001", "010", "011", '0', '-', "00"), -- i=4248
      ("1010101100010010", '1', '1', "10", "001", "010", "011", '0', '-', "00"), -- i=4249
      ("1010101100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4250
      ("1011001100010010", '0', '1', "11", "001", "010", "011", '0', '-', "00"), -- i=4251
      ("1011101100010010", '1', '1', "11", "001", "010", "011", '0', '-', "00"), -- i=4252
      ("1011101100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4253
      ("0101001100010000", '0', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4254
      ("0101101100010000", '1', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4255
      ("0101101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4256
      ("0100001100010000", '0', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4257
      ("0100101100010000", '1', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4258
      ("0100101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4259
      ("0000001101100000", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4260
      ("0000101101100000", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4261
      ("0000101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4262
      ("1000001100010011", '0', '1', "00", "001", "011", "011", '0', '-', "00"), -- i=4263
      ("1000101100010011", '1', '1', "00", "001", "011", "011", '0', '-', "00"), -- i=4264
      ("1000101100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4265
      ("1001001100010011", '0', '1', "01", "001", "011", "011", '0', '-', "00"), -- i=4266
      ("1001101100010011", '1', '1', "01", "001", "011", "011", '0', '-', "00"), -- i=4267
      ("1001101100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4268
      ("1010001100010011", '0', '1', "10", "001", "011", "011", '0', '-', "00"), -- i=4269
      ("1010101100010011", '1', '1', "10", "001", "011", "011", '0', '-', "00"), -- i=4270
      ("1010101100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4271
      ("1011001100010011", '0', '1', "11", "001", "011", "011", '0', '-', "00"), -- i=4272
      ("1011101100010011", '1', '1', "11", "001", "011", "011", '0', '-', "00"), -- i=4273
      ("1011101100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4274
      ("0101001100010000", '0', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4275
      ("0101101100010000", '1', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4276
      ("0101101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4277
      ("0100001100010000", '0', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4278
      ("0100101100010000", '1', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4279
      ("0100101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4280
      ("0000001101010110", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4281
      ("0000101101010110", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4282
      ("0000101101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4283
      ("1000001100010100", '0', '1', "00", "001", "100", "011", '0', '-', "00"), -- i=4284
      ("1000101100010100", '1', '1', "00", "001", "100", "011", '0', '-', "00"), -- i=4285
      ("1000101100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4286
      ("1001001100010100", '0', '1', "01", "001", "100", "011", '0', '-', "00"), -- i=4287
      ("1001101100010100", '1', '1', "01", "001", "100", "011", '0', '-', "00"), -- i=4288
      ("1001101100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4289
      ("1010001100010100", '0', '1', "10", "001", "100", "011", '0', '-', "00"), -- i=4290
      ("1010101100010100", '1', '1', "10", "001", "100", "011", '0', '-', "00"), -- i=4291
      ("1010101100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4292
      ("1011001100010100", '0', '1', "11", "001", "100", "011", '0', '-', "00"), -- i=4293
      ("1011101100010100", '1', '1', "11", "001", "100", "011", '0', '-', "00"), -- i=4294
      ("1011101100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4295
      ("0101001100010000", '0', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4296
      ("0101101100010000", '1', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4297
      ("0101101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4298
      ("0100001100010000", '0', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4299
      ("0100101100010000", '1', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4300
      ("0100101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4301
      ("0000001101111001", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4302
      ("0000101101111001", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4303
      ("0000101101111001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4304
      ("1000001100010101", '0', '1', "00", "001", "101", "011", '0', '-', "00"), -- i=4305
      ("1000101100010101", '1', '1', "00", "001", "101", "011", '0', '-', "00"), -- i=4306
      ("1000101100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4307
      ("1001001100010101", '0', '1', "01", "001", "101", "011", '0', '-', "00"), -- i=4308
      ("1001101100010101", '1', '1', "01", "001", "101", "011", '0', '-', "00"), -- i=4309
      ("1001101100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4310
      ("1010001100010101", '0', '1', "10", "001", "101", "011", '0', '-', "00"), -- i=4311
      ("1010101100010101", '1', '1', "10", "001", "101", "011", '0', '-', "00"), -- i=4312
      ("1010101100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4313
      ("1011001100010101", '0', '1', "11", "001", "101", "011", '0', '-', "00"), -- i=4314
      ("1011101100010101", '1', '1', "11", "001", "101", "011", '0', '-', "00"), -- i=4315
      ("1011101100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4316
      ("0101001100010000", '0', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4317
      ("0101101100010000", '1', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4318
      ("0101101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4319
      ("0100001100010000", '0', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4320
      ("0100101100010000", '1', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4321
      ("0100101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4322
      ("0000001110101100", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4323
      ("0000101110101100", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4324
      ("0000101110101100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4325
      ("1000001100010110", '0', '1', "00", "001", "110", "011", '0', '-', "00"), -- i=4326
      ("1000101100010110", '1', '1', "00", "001", "110", "011", '0', '-', "00"), -- i=4327
      ("1000101100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4328
      ("1001001100010110", '0', '1', "01", "001", "110", "011", '0', '-', "00"), -- i=4329
      ("1001101100010110", '1', '1', "01", "001", "110", "011", '0', '-', "00"), -- i=4330
      ("1001101100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4331
      ("1010001100010110", '0', '1', "10", "001", "110", "011", '0', '-', "00"), -- i=4332
      ("1010101100010110", '1', '1', "10", "001", "110", "011", '0', '-', "00"), -- i=4333
      ("1010101100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4334
      ("1011001100010110", '0', '1', "11", "001", "110", "011", '0', '-', "00"), -- i=4335
      ("1011101100010110", '1', '1', "11", "001", "110", "011", '0', '-', "00"), -- i=4336
      ("1011101100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4337
      ("0101001100010000", '0', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4338
      ("0101101100010000", '1', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4339
      ("0101101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4340
      ("0100001100010000", '0', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4341
      ("0100101100010000", '1', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4342
      ("0100101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4343
      ("0000001111000100", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4344
      ("0000101111000100", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4345
      ("0000101111000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4346
      ("1000001100010111", '0', '1', "00", "001", "111", "011", '0', '-', "00"), -- i=4347
      ("1000101100010111", '1', '1', "00", "001", "111", "011", '0', '-', "00"), -- i=4348
      ("1000101100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4349
      ("1001001100010111", '0', '1', "01", "001", "111", "011", '0', '-', "00"), -- i=4350
      ("1001101100010111", '1', '1', "01", "001", "111", "011", '0', '-', "00"), -- i=4351
      ("1001101100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4352
      ("1010001100010111", '0', '1', "10", "001", "111", "011", '0', '-', "00"), -- i=4353
      ("1010101100010111", '1', '1', "10", "001", "111", "011", '0', '-', "00"), -- i=4354
      ("1010101100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4355
      ("1011001100010111", '0', '1', "11", "001", "111", "011", '0', '-', "00"), -- i=4356
      ("1011101100010111", '1', '1', "11", "001", "111", "011", '0', '-', "00"), -- i=4357
      ("1011101100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4358
      ("0101001100010000", '0', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4359
      ("0101101100010000", '1', '1', "--", "001", "---", "011", '0', '1', "01"), -- i=4360
      ("0101101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4361
      ("0100001100010000", '0', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4362
      ("0100101100010000", '1', '0', "--", "001", "011", "---", '1', '-', "--"), -- i=4363
      ("0100101100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4364
      ("0000001101111010", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4365
      ("0000101101111010", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4366
      ("0000101101111010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4367
      ("1000001100100000", '0', '1', "00", "010", "000", "011", '0', '-', "00"), -- i=4368
      ("1000101100100000", '1', '1', "00", "010", "000", "011", '0', '-', "00"), -- i=4369
      ("1000101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4370
      ("1001001100100000", '0', '1', "01", "010", "000", "011", '0', '-', "00"), -- i=4371
      ("1001101100100000", '1', '1', "01", "010", "000", "011", '0', '-', "00"), -- i=4372
      ("1001101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4373
      ("1010001100100000", '0', '1', "10", "010", "000", "011", '0', '-', "00"), -- i=4374
      ("1010101100100000", '1', '1', "10", "010", "000", "011", '0', '-', "00"), -- i=4375
      ("1010101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4376
      ("1011001100100000", '0', '1', "11", "010", "000", "011", '0', '-', "00"), -- i=4377
      ("1011101100100000", '1', '1', "11", "010", "000", "011", '0', '-', "00"), -- i=4378
      ("1011101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4379
      ("0101001100100000", '0', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4380
      ("0101101100100000", '1', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4381
      ("0101101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4382
      ("0100001100100000", '0', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4383
      ("0100101100100000", '1', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4384
      ("0100101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4385
      ("0000001100000101", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4386
      ("0000101100000101", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4387
      ("0000101100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4388
      ("1000001100100001", '0', '1', "00", "010", "001", "011", '0', '-', "00"), -- i=4389
      ("1000101100100001", '1', '1', "00", "010", "001", "011", '0', '-', "00"), -- i=4390
      ("1000101100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4391
      ("1001001100100001", '0', '1', "01", "010", "001", "011", '0', '-', "00"), -- i=4392
      ("1001101100100001", '1', '1', "01", "010", "001", "011", '0', '-', "00"), -- i=4393
      ("1001101100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4394
      ("1010001100100001", '0', '1', "10", "010", "001", "011", '0', '-', "00"), -- i=4395
      ("1010101100100001", '1', '1', "10", "010", "001", "011", '0', '-', "00"), -- i=4396
      ("1010101100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4397
      ("1011001100100001", '0', '1', "11", "010", "001", "011", '0', '-', "00"), -- i=4398
      ("1011101100100001", '1', '1', "11", "010", "001", "011", '0', '-', "00"), -- i=4399
      ("1011101100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4400
      ("0101001100100000", '0', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4401
      ("0101101100100000", '1', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4402
      ("0101101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4403
      ("0100001100100000", '0', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4404
      ("0100101100100000", '1', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4405
      ("0100101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4406
      ("0000001110111110", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4407
      ("0000101110111110", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4408
      ("0000101110111110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4409
      ("1000001100100010", '0', '1', "00", "010", "010", "011", '0', '-', "00"), -- i=4410
      ("1000101100100010", '1', '1', "00", "010", "010", "011", '0', '-', "00"), -- i=4411
      ("1000101100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4412
      ("1001001100100010", '0', '1', "01", "010", "010", "011", '0', '-', "00"), -- i=4413
      ("1001101100100010", '1', '1', "01", "010", "010", "011", '0', '-', "00"), -- i=4414
      ("1001101100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4415
      ("1010001100100010", '0', '1', "10", "010", "010", "011", '0', '-', "00"), -- i=4416
      ("1010101100100010", '1', '1', "10", "010", "010", "011", '0', '-', "00"), -- i=4417
      ("1010101100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4418
      ("1011001100100010", '0', '1', "11", "010", "010", "011", '0', '-', "00"), -- i=4419
      ("1011101100100010", '1', '1', "11", "010", "010", "011", '0', '-', "00"), -- i=4420
      ("1011101100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4421
      ("0101001100100000", '0', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4422
      ("0101101100100000", '1', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4423
      ("0101101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4424
      ("0100001100100000", '0', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4425
      ("0100101100100000", '1', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4426
      ("0100101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4427
      ("0000001100100000", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4428
      ("0000101100100000", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4429
      ("0000101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4430
      ("1000001100100011", '0', '1', "00", "010", "011", "011", '0', '-', "00"), -- i=4431
      ("1000101100100011", '1', '1', "00", "010", "011", "011", '0', '-', "00"), -- i=4432
      ("1000101100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4433
      ("1001001100100011", '0', '1', "01", "010", "011", "011", '0', '-', "00"), -- i=4434
      ("1001101100100011", '1', '1', "01", "010", "011", "011", '0', '-', "00"), -- i=4435
      ("1001101100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4436
      ("1010001100100011", '0', '1', "10", "010", "011", "011", '0', '-', "00"), -- i=4437
      ("1010101100100011", '1', '1', "10", "010", "011", "011", '0', '-', "00"), -- i=4438
      ("1010101100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4439
      ("1011001100100011", '0', '1', "11", "010", "011", "011", '0', '-', "00"), -- i=4440
      ("1011101100100011", '1', '1', "11", "010", "011", "011", '0', '-', "00"), -- i=4441
      ("1011101100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4442
      ("0101001100100000", '0', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4443
      ("0101101100100000", '1', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4444
      ("0101101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4445
      ("0100001100100000", '0', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4446
      ("0100101100100000", '1', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4447
      ("0100101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4448
      ("0000001111100100", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4449
      ("0000101111100100", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4450
      ("0000101111100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4451
      ("1000001100100100", '0', '1', "00", "010", "100", "011", '0', '-', "00"), -- i=4452
      ("1000101100100100", '1', '1', "00", "010", "100", "011", '0', '-', "00"), -- i=4453
      ("1000101100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4454
      ("1001001100100100", '0', '1', "01", "010", "100", "011", '0', '-', "00"), -- i=4455
      ("1001101100100100", '1', '1', "01", "010", "100", "011", '0', '-', "00"), -- i=4456
      ("1001101100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4457
      ("1010001100100100", '0', '1', "10", "010", "100", "011", '0', '-', "00"), -- i=4458
      ("1010101100100100", '1', '1', "10", "010", "100", "011", '0', '-', "00"), -- i=4459
      ("1010101100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4460
      ("1011001100100100", '0', '1', "11", "010", "100", "011", '0', '-', "00"), -- i=4461
      ("1011101100100100", '1', '1', "11", "010", "100", "011", '0', '-', "00"), -- i=4462
      ("1011101100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4463
      ("0101001100100000", '0', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4464
      ("0101101100100000", '1', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4465
      ("0101101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4466
      ("0100001100100000", '0', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4467
      ("0100101100100000", '1', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4468
      ("0100101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4469
      ("0000001100100010", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4470
      ("0000101100100010", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4471
      ("0000101100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4472
      ("1000001100100101", '0', '1', "00", "010", "101", "011", '0', '-', "00"), -- i=4473
      ("1000101100100101", '1', '1', "00", "010", "101", "011", '0', '-', "00"), -- i=4474
      ("1000101100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4475
      ("1001001100100101", '0', '1', "01", "010", "101", "011", '0', '-', "00"), -- i=4476
      ("1001101100100101", '1', '1', "01", "010", "101", "011", '0', '-', "00"), -- i=4477
      ("1001101100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4478
      ("1010001100100101", '0', '1', "10", "010", "101", "011", '0', '-', "00"), -- i=4479
      ("1010101100100101", '1', '1', "10", "010", "101", "011", '0', '-', "00"), -- i=4480
      ("1010101100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4481
      ("1011001100100101", '0', '1', "11", "010", "101", "011", '0', '-', "00"), -- i=4482
      ("1011101100100101", '1', '1', "11", "010", "101", "011", '0', '-', "00"), -- i=4483
      ("1011101100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4484
      ("0101001100100000", '0', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4485
      ("0101101100100000", '1', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4486
      ("0101101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4487
      ("0100001100100000", '0', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4488
      ("0100101100100000", '1', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4489
      ("0100101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4490
      ("0000001100101101", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4491
      ("0000101100101101", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4492
      ("0000101100101101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4493
      ("1000001100100110", '0', '1', "00", "010", "110", "011", '0', '-', "00"), -- i=4494
      ("1000101100100110", '1', '1', "00", "010", "110", "011", '0', '-', "00"), -- i=4495
      ("1000101100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4496
      ("1001001100100110", '0', '1', "01", "010", "110", "011", '0', '-', "00"), -- i=4497
      ("1001101100100110", '1', '1', "01", "010", "110", "011", '0', '-', "00"), -- i=4498
      ("1001101100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4499
      ("1010001100100110", '0', '1', "10", "010", "110", "011", '0', '-', "00"), -- i=4500
      ("1010101100100110", '1', '1', "10", "010", "110", "011", '0', '-', "00"), -- i=4501
      ("1010101100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4502
      ("1011001100100110", '0', '1', "11", "010", "110", "011", '0', '-', "00"), -- i=4503
      ("1011101100100110", '1', '1', "11", "010", "110", "011", '0', '-', "00"), -- i=4504
      ("1011101100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4505
      ("0101001100100000", '0', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4506
      ("0101101100100000", '1', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4507
      ("0101101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4508
      ("0100001100100000", '0', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4509
      ("0100101100100000", '1', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4510
      ("0100101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4511
      ("0000001100000001", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4512
      ("0000101100000001", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4513
      ("0000101100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4514
      ("1000001100100111", '0', '1', "00", "010", "111", "011", '0', '-', "00"), -- i=4515
      ("1000101100100111", '1', '1', "00", "010", "111", "011", '0', '-', "00"), -- i=4516
      ("1000101100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4517
      ("1001001100100111", '0', '1', "01", "010", "111", "011", '0', '-', "00"), -- i=4518
      ("1001101100100111", '1', '1', "01", "010", "111", "011", '0', '-', "00"), -- i=4519
      ("1001101100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4520
      ("1010001100100111", '0', '1', "10", "010", "111", "011", '0', '-', "00"), -- i=4521
      ("1010101100100111", '1', '1', "10", "010", "111", "011", '0', '-', "00"), -- i=4522
      ("1010101100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4523
      ("1011001100100111", '0', '1', "11", "010", "111", "011", '0', '-', "00"), -- i=4524
      ("1011101100100111", '1', '1', "11", "010", "111", "011", '0', '-', "00"), -- i=4525
      ("1011101100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4526
      ("0101001100100000", '0', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4527
      ("0101101100100000", '1', '1', "--", "010", "---", "011", '0', '1', "01"), -- i=4528
      ("0101101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4529
      ("0100001100100000", '0', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4530
      ("0100101100100000", '1', '0', "--", "010", "011", "---", '1', '-', "--"), -- i=4531
      ("0100101100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4532
      ("0000001100011010", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4533
      ("0000101100011010", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4534
      ("0000101100011010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4535
      ("1000001100110000", '0', '1', "00", "011", "000", "011", '0', '-', "00"), -- i=4536
      ("1000101100110000", '1', '1', "00", "011", "000", "011", '0', '-', "00"), -- i=4537
      ("1000101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4538
      ("1001001100110000", '0', '1', "01", "011", "000", "011", '0', '-', "00"), -- i=4539
      ("1001101100110000", '1', '1', "01", "011", "000", "011", '0', '-', "00"), -- i=4540
      ("1001101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4541
      ("1010001100110000", '0', '1', "10", "011", "000", "011", '0', '-', "00"), -- i=4542
      ("1010101100110000", '1', '1', "10", "011", "000", "011", '0', '-', "00"), -- i=4543
      ("1010101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4544
      ("1011001100110000", '0', '1', "11", "011", "000", "011", '0', '-', "00"), -- i=4545
      ("1011101100110000", '1', '1', "11", "011", "000", "011", '0', '-', "00"), -- i=4546
      ("1011101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4547
      ("0101001100110000", '0', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4548
      ("0101101100110000", '1', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4549
      ("0101101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4550
      ("0100001100110000", '0', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4551
      ("0100101100110000", '1', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4552
      ("0100101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4553
      ("0000001110100111", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4554
      ("0000101110100111", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4555
      ("0000101110100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4556
      ("1000001100110001", '0', '1', "00", "011", "001", "011", '0', '-', "00"), -- i=4557
      ("1000101100110001", '1', '1', "00", "011", "001", "011", '0', '-', "00"), -- i=4558
      ("1000101100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4559
      ("1001001100110001", '0', '1', "01", "011", "001", "011", '0', '-', "00"), -- i=4560
      ("1001101100110001", '1', '1', "01", "011", "001", "011", '0', '-', "00"), -- i=4561
      ("1001101100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4562
      ("1010001100110001", '0', '1', "10", "011", "001", "011", '0', '-', "00"), -- i=4563
      ("1010101100110001", '1', '1', "10", "011", "001", "011", '0', '-', "00"), -- i=4564
      ("1010101100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4565
      ("1011001100110001", '0', '1', "11", "011", "001", "011", '0', '-', "00"), -- i=4566
      ("1011101100110001", '1', '1', "11", "011", "001", "011", '0', '-', "00"), -- i=4567
      ("1011101100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4568
      ("0101001100110000", '0', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4569
      ("0101101100110000", '1', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4570
      ("0101101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4571
      ("0100001100110000", '0', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4572
      ("0100101100110000", '1', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4573
      ("0100101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4574
      ("0000001110110111", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4575
      ("0000101110110111", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4576
      ("0000101110110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4577
      ("1000001100110010", '0', '1', "00", "011", "010", "011", '0', '-', "00"), -- i=4578
      ("1000101100110010", '1', '1', "00", "011", "010", "011", '0', '-', "00"), -- i=4579
      ("1000101100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4580
      ("1001001100110010", '0', '1', "01", "011", "010", "011", '0', '-', "00"), -- i=4581
      ("1001101100110010", '1', '1', "01", "011", "010", "011", '0', '-', "00"), -- i=4582
      ("1001101100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4583
      ("1010001100110010", '0', '1', "10", "011", "010", "011", '0', '-', "00"), -- i=4584
      ("1010101100110010", '1', '1', "10", "011", "010", "011", '0', '-', "00"), -- i=4585
      ("1010101100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4586
      ("1011001100110010", '0', '1', "11", "011", "010", "011", '0', '-', "00"), -- i=4587
      ("1011101100110010", '1', '1', "11", "011", "010", "011", '0', '-', "00"), -- i=4588
      ("1011101100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4589
      ("0101001100110000", '0', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4590
      ("0101101100110000", '1', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4591
      ("0101101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4592
      ("0100001100110000", '0', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4593
      ("0100101100110000", '1', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4594
      ("0100101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4595
      ("0000001100101000", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4596
      ("0000101100101000", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4597
      ("0000101100101000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4598
      ("1000001100110011", '0', '1', "00", "011", "011", "011", '0', '-', "00"), -- i=4599
      ("1000101100110011", '1', '1', "00", "011", "011", "011", '0', '-', "00"), -- i=4600
      ("1000101100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4601
      ("1001001100110011", '0', '1', "01", "011", "011", "011", '0', '-', "00"), -- i=4602
      ("1001101100110011", '1', '1', "01", "011", "011", "011", '0', '-', "00"), -- i=4603
      ("1001101100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4604
      ("1010001100110011", '0', '1', "10", "011", "011", "011", '0', '-', "00"), -- i=4605
      ("1010101100110011", '1', '1', "10", "011", "011", "011", '0', '-', "00"), -- i=4606
      ("1010101100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4607
      ("1011001100110011", '0', '1', "11", "011", "011", "011", '0', '-', "00"), -- i=4608
      ("1011101100110011", '1', '1', "11", "011", "011", "011", '0', '-', "00"), -- i=4609
      ("1011101100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4610
      ("0101001100110000", '0', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4611
      ("0101101100110000", '1', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4612
      ("0101101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4613
      ("0100001100110000", '0', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4614
      ("0100101100110000", '1', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4615
      ("0100101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4616
      ("0000001100000010", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4617
      ("0000101100000010", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4618
      ("0000101100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4619
      ("1000001100110100", '0', '1', "00", "011", "100", "011", '0', '-', "00"), -- i=4620
      ("1000101100110100", '1', '1', "00", "011", "100", "011", '0', '-', "00"), -- i=4621
      ("1000101100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4622
      ("1001001100110100", '0', '1', "01", "011", "100", "011", '0', '-', "00"), -- i=4623
      ("1001101100110100", '1', '1', "01", "011", "100", "011", '0', '-', "00"), -- i=4624
      ("1001101100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4625
      ("1010001100110100", '0', '1', "10", "011", "100", "011", '0', '-', "00"), -- i=4626
      ("1010101100110100", '1', '1', "10", "011", "100", "011", '0', '-', "00"), -- i=4627
      ("1010101100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4628
      ("1011001100110100", '0', '1', "11", "011", "100", "011", '0', '-', "00"), -- i=4629
      ("1011101100110100", '1', '1', "11", "011", "100", "011", '0', '-', "00"), -- i=4630
      ("1011101100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4631
      ("0101001100110000", '0', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4632
      ("0101101100110000", '1', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4633
      ("0101101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4634
      ("0100001100110000", '0', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4635
      ("0100101100110000", '1', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4636
      ("0100101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4637
      ("0000001110100111", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4638
      ("0000101110100111", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4639
      ("0000101110100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4640
      ("1000001100110101", '0', '1', "00", "011", "101", "011", '0', '-', "00"), -- i=4641
      ("1000101100110101", '1', '1', "00", "011", "101", "011", '0', '-', "00"), -- i=4642
      ("1000101100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4643
      ("1001001100110101", '0', '1', "01", "011", "101", "011", '0', '-', "00"), -- i=4644
      ("1001101100110101", '1', '1', "01", "011", "101", "011", '0', '-', "00"), -- i=4645
      ("1001101100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4646
      ("1010001100110101", '0', '1', "10", "011", "101", "011", '0', '-', "00"), -- i=4647
      ("1010101100110101", '1', '1', "10", "011", "101", "011", '0', '-', "00"), -- i=4648
      ("1010101100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4649
      ("1011001100110101", '0', '1', "11", "011", "101", "011", '0', '-', "00"), -- i=4650
      ("1011101100110101", '1', '1', "11", "011", "101", "011", '0', '-', "00"), -- i=4651
      ("1011101100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4652
      ("0101001100110000", '0', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4653
      ("0101101100110000", '1', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4654
      ("0101101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4655
      ("0100001100110000", '0', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4656
      ("0100101100110000", '1', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4657
      ("0100101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4658
      ("0000001110010100", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4659
      ("0000101110010100", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4660
      ("0000101110010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4661
      ("1000001100110110", '0', '1', "00", "011", "110", "011", '0', '-', "00"), -- i=4662
      ("1000101100110110", '1', '1', "00", "011", "110", "011", '0', '-', "00"), -- i=4663
      ("1000101100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4664
      ("1001001100110110", '0', '1', "01", "011", "110", "011", '0', '-', "00"), -- i=4665
      ("1001101100110110", '1', '1', "01", "011", "110", "011", '0', '-', "00"), -- i=4666
      ("1001101100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4667
      ("1010001100110110", '0', '1', "10", "011", "110", "011", '0', '-', "00"), -- i=4668
      ("1010101100110110", '1', '1', "10", "011", "110", "011", '0', '-', "00"), -- i=4669
      ("1010101100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4670
      ("1011001100110110", '0', '1', "11", "011", "110", "011", '0', '-', "00"), -- i=4671
      ("1011101100110110", '1', '1', "11", "011", "110", "011", '0', '-', "00"), -- i=4672
      ("1011101100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4673
      ("0101001100110000", '0', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4674
      ("0101101100110000", '1', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4675
      ("0101101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4676
      ("0100001100110000", '0', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4677
      ("0100101100110000", '1', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4678
      ("0100101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4679
      ("0000001100110111", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4680
      ("0000101100110111", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4681
      ("0000101100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4682
      ("1000001100110111", '0', '1', "00", "011", "111", "011", '0', '-', "00"), -- i=4683
      ("1000101100110111", '1', '1', "00", "011", "111", "011", '0', '-', "00"), -- i=4684
      ("1000101100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4685
      ("1001001100110111", '0', '1', "01", "011", "111", "011", '0', '-', "00"), -- i=4686
      ("1001101100110111", '1', '1', "01", "011", "111", "011", '0', '-', "00"), -- i=4687
      ("1001101100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4688
      ("1010001100110111", '0', '1', "10", "011", "111", "011", '0', '-', "00"), -- i=4689
      ("1010101100110111", '1', '1', "10", "011", "111", "011", '0', '-', "00"), -- i=4690
      ("1010101100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4691
      ("1011001100110111", '0', '1', "11", "011", "111", "011", '0', '-', "00"), -- i=4692
      ("1011101100110111", '1', '1', "11", "011", "111", "011", '0', '-', "00"), -- i=4693
      ("1011101100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4694
      ("0101001100110000", '0', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4695
      ("0101101100110000", '1', '1', "--", "011", "---", "011", '0', '1', "01"), -- i=4696
      ("0101101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4697
      ("0100001100110000", '0', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4698
      ("0100101100110000", '1', '0', "--", "011", "011", "---", '1', '-', "--"), -- i=4699
      ("0100101100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4700
      ("0000001111000100", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4701
      ("0000101111000100", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4702
      ("0000101111000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4703
      ("1000001101000000", '0', '1', "00", "100", "000", "011", '0', '-', "00"), -- i=4704
      ("1000101101000000", '1', '1', "00", "100", "000", "011", '0', '-', "00"), -- i=4705
      ("1000101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4706
      ("1001001101000000", '0', '1', "01", "100", "000", "011", '0', '-', "00"), -- i=4707
      ("1001101101000000", '1', '1', "01", "100", "000", "011", '0', '-', "00"), -- i=4708
      ("1001101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4709
      ("1010001101000000", '0', '1', "10", "100", "000", "011", '0', '-', "00"), -- i=4710
      ("1010101101000000", '1', '1', "10", "100", "000", "011", '0', '-', "00"), -- i=4711
      ("1010101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4712
      ("1011001101000000", '0', '1', "11", "100", "000", "011", '0', '-', "00"), -- i=4713
      ("1011101101000000", '1', '1', "11", "100", "000", "011", '0', '-', "00"), -- i=4714
      ("1011101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4715
      ("0101001101000000", '0', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4716
      ("0101101101000000", '1', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4717
      ("0101101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4718
      ("0100001101000000", '0', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4719
      ("0100101101000000", '1', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4720
      ("0100101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4721
      ("0000001100001101", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4722
      ("0000101100001101", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4723
      ("0000101100001101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4724
      ("1000001101000001", '0', '1', "00", "100", "001", "011", '0', '-', "00"), -- i=4725
      ("1000101101000001", '1', '1', "00", "100", "001", "011", '0', '-', "00"), -- i=4726
      ("1000101101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4727
      ("1001001101000001", '0', '1', "01", "100", "001", "011", '0', '-', "00"), -- i=4728
      ("1001101101000001", '1', '1', "01", "100", "001", "011", '0', '-', "00"), -- i=4729
      ("1001101101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4730
      ("1010001101000001", '0', '1', "10", "100", "001", "011", '0', '-', "00"), -- i=4731
      ("1010101101000001", '1', '1', "10", "100", "001", "011", '0', '-', "00"), -- i=4732
      ("1010101101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4733
      ("1011001101000001", '0', '1', "11", "100", "001", "011", '0', '-', "00"), -- i=4734
      ("1011101101000001", '1', '1', "11", "100", "001", "011", '0', '-', "00"), -- i=4735
      ("1011101101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4736
      ("0101001101000000", '0', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4737
      ("0101101101000000", '1', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4738
      ("0101101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4739
      ("0100001101000000", '0', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4740
      ("0100101101000000", '1', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4741
      ("0100101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4742
      ("0000001100011000", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4743
      ("0000101100011000", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4744
      ("0000101100011000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4745
      ("1000001101000010", '0', '1', "00", "100", "010", "011", '0', '-', "00"), -- i=4746
      ("1000101101000010", '1', '1', "00", "100", "010", "011", '0', '-', "00"), -- i=4747
      ("1000101101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4748
      ("1001001101000010", '0', '1', "01", "100", "010", "011", '0', '-', "00"), -- i=4749
      ("1001101101000010", '1', '1', "01", "100", "010", "011", '0', '-', "00"), -- i=4750
      ("1001101101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4751
      ("1010001101000010", '0', '1', "10", "100", "010", "011", '0', '-', "00"), -- i=4752
      ("1010101101000010", '1', '1', "10", "100", "010", "011", '0', '-', "00"), -- i=4753
      ("1010101101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4754
      ("1011001101000010", '0', '1', "11", "100", "010", "011", '0', '-', "00"), -- i=4755
      ("1011101101000010", '1', '1', "11", "100", "010", "011", '0', '-', "00"), -- i=4756
      ("1011101101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4757
      ("0101001101000000", '0', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4758
      ("0101101101000000", '1', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4759
      ("0101101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4760
      ("0100001101000000", '0', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4761
      ("0100101101000000", '1', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4762
      ("0100101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4763
      ("0000001110101111", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4764
      ("0000101110101111", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4765
      ("0000101110101111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4766
      ("1000001101000011", '0', '1', "00", "100", "011", "011", '0', '-', "00"), -- i=4767
      ("1000101101000011", '1', '1', "00", "100", "011", "011", '0', '-', "00"), -- i=4768
      ("1000101101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4769
      ("1001001101000011", '0', '1', "01", "100", "011", "011", '0', '-', "00"), -- i=4770
      ("1001101101000011", '1', '1', "01", "100", "011", "011", '0', '-', "00"), -- i=4771
      ("1001101101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4772
      ("1010001101000011", '0', '1', "10", "100", "011", "011", '0', '-', "00"), -- i=4773
      ("1010101101000011", '1', '1', "10", "100", "011", "011", '0', '-', "00"), -- i=4774
      ("1010101101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4775
      ("1011001101000011", '0', '1', "11", "100", "011", "011", '0', '-', "00"), -- i=4776
      ("1011101101000011", '1', '1', "11", "100", "011", "011", '0', '-', "00"), -- i=4777
      ("1011101101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4778
      ("0101001101000000", '0', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4779
      ("0101101101000000", '1', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4780
      ("0101101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4781
      ("0100001101000000", '0', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4782
      ("0100101101000000", '1', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4783
      ("0100101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4784
      ("0000001110000001", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4785
      ("0000101110000001", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4786
      ("0000101110000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4787
      ("1000001101000100", '0', '1', "00", "100", "100", "011", '0', '-', "00"), -- i=4788
      ("1000101101000100", '1', '1', "00", "100", "100", "011", '0', '-', "00"), -- i=4789
      ("1000101101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4790
      ("1001001101000100", '0', '1', "01", "100", "100", "011", '0', '-', "00"), -- i=4791
      ("1001101101000100", '1', '1', "01", "100", "100", "011", '0', '-', "00"), -- i=4792
      ("1001101101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4793
      ("1010001101000100", '0', '1', "10", "100", "100", "011", '0', '-', "00"), -- i=4794
      ("1010101101000100", '1', '1', "10", "100", "100", "011", '0', '-', "00"), -- i=4795
      ("1010101101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4796
      ("1011001101000100", '0', '1', "11", "100", "100", "011", '0', '-', "00"), -- i=4797
      ("1011101101000100", '1', '1', "11", "100", "100", "011", '0', '-', "00"), -- i=4798
      ("1011101101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4799
      ("0101001101000000", '0', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4800
      ("0101101101000000", '1', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4801
      ("0101101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4802
      ("0100001101000000", '0', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4803
      ("0100101101000000", '1', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4804
      ("0100101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4805
      ("0000001101100011", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4806
      ("0000101101100011", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4807
      ("0000101101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4808
      ("1000001101000101", '0', '1', "00", "100", "101", "011", '0', '-', "00"), -- i=4809
      ("1000101101000101", '1', '1', "00", "100", "101", "011", '0', '-', "00"), -- i=4810
      ("1000101101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4811
      ("1001001101000101", '0', '1', "01", "100", "101", "011", '0', '-', "00"), -- i=4812
      ("1001101101000101", '1', '1', "01", "100", "101", "011", '0', '-', "00"), -- i=4813
      ("1001101101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4814
      ("1010001101000101", '0', '1', "10", "100", "101", "011", '0', '-', "00"), -- i=4815
      ("1010101101000101", '1', '1', "10", "100", "101", "011", '0', '-', "00"), -- i=4816
      ("1010101101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4817
      ("1011001101000101", '0', '1', "11", "100", "101", "011", '0', '-', "00"), -- i=4818
      ("1011101101000101", '1', '1', "11", "100", "101", "011", '0', '-', "00"), -- i=4819
      ("1011101101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4820
      ("0101001101000000", '0', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4821
      ("0101101101000000", '1', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4822
      ("0101101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4823
      ("0100001101000000", '0', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4824
      ("0100101101000000", '1', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4825
      ("0100101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4826
      ("0000001111010110", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4827
      ("0000101111010110", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4828
      ("0000101111010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4829
      ("1000001101000110", '0', '1', "00", "100", "110", "011", '0', '-', "00"), -- i=4830
      ("1000101101000110", '1', '1', "00", "100", "110", "011", '0', '-', "00"), -- i=4831
      ("1000101101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4832
      ("1001001101000110", '0', '1', "01", "100", "110", "011", '0', '-', "00"), -- i=4833
      ("1001101101000110", '1', '1', "01", "100", "110", "011", '0', '-', "00"), -- i=4834
      ("1001101101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4835
      ("1010001101000110", '0', '1', "10", "100", "110", "011", '0', '-', "00"), -- i=4836
      ("1010101101000110", '1', '1', "10", "100", "110", "011", '0', '-', "00"), -- i=4837
      ("1010101101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4838
      ("1011001101000110", '0', '1', "11", "100", "110", "011", '0', '-', "00"), -- i=4839
      ("1011101101000110", '1', '1', "11", "100", "110", "011", '0', '-', "00"), -- i=4840
      ("1011101101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4841
      ("0101001101000000", '0', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4842
      ("0101101101000000", '1', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4843
      ("0101101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4844
      ("0100001101000000", '0', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4845
      ("0100101101000000", '1', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4846
      ("0100101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4847
      ("0000001100010001", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4848
      ("0000101100010001", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4849
      ("0000101100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4850
      ("1000001101000111", '0', '1', "00", "100", "111", "011", '0', '-', "00"), -- i=4851
      ("1000101101000111", '1', '1', "00", "100", "111", "011", '0', '-', "00"), -- i=4852
      ("1000101101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4853
      ("1001001101000111", '0', '1', "01", "100", "111", "011", '0', '-', "00"), -- i=4854
      ("1001101101000111", '1', '1', "01", "100", "111", "011", '0', '-', "00"), -- i=4855
      ("1001101101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4856
      ("1010001101000111", '0', '1', "10", "100", "111", "011", '0', '-', "00"), -- i=4857
      ("1010101101000111", '1', '1', "10", "100", "111", "011", '0', '-', "00"), -- i=4858
      ("1010101101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4859
      ("1011001101000111", '0', '1', "11", "100", "111", "011", '0', '-', "00"), -- i=4860
      ("1011101101000111", '1', '1', "11", "100", "111", "011", '0', '-', "00"), -- i=4861
      ("1011101101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4862
      ("0101001101000000", '0', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4863
      ("0101101101000000", '1', '1', "--", "100", "---", "011", '0', '1', "01"), -- i=4864
      ("0101101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4865
      ("0100001101000000", '0', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4866
      ("0100101101000000", '1', '0', "--", "100", "011", "---", '1', '-', "--"), -- i=4867
      ("0100101101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4868
      ("0000001100110101", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4869
      ("0000101100110101", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4870
      ("0000101100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4871
      ("1000001101010000", '0', '1', "00", "101", "000", "011", '0', '-', "00"), -- i=4872
      ("1000101101010000", '1', '1', "00", "101", "000", "011", '0', '-', "00"), -- i=4873
      ("1000101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4874
      ("1001001101010000", '0', '1', "01", "101", "000", "011", '0', '-', "00"), -- i=4875
      ("1001101101010000", '1', '1', "01", "101", "000", "011", '0', '-', "00"), -- i=4876
      ("1001101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4877
      ("1010001101010000", '0', '1', "10", "101", "000", "011", '0', '-', "00"), -- i=4878
      ("1010101101010000", '1', '1', "10", "101", "000", "011", '0', '-', "00"), -- i=4879
      ("1010101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4880
      ("1011001101010000", '0', '1', "11", "101", "000", "011", '0', '-', "00"), -- i=4881
      ("1011101101010000", '1', '1', "11", "101", "000", "011", '0', '-', "00"), -- i=4882
      ("1011101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4883
      ("0101001101010000", '0', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=4884
      ("0101101101010000", '1', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=4885
      ("0101101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4886
      ("0100001101010000", '0', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=4887
      ("0100101101010000", '1', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=4888
      ("0100101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4889
      ("0000001101110001", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4890
      ("0000101101110001", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4891
      ("0000101101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4892
      ("1000001101010001", '0', '1', "00", "101", "001", "011", '0', '-', "00"), -- i=4893
      ("1000101101010001", '1', '1', "00", "101", "001", "011", '0', '-', "00"), -- i=4894
      ("1000101101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4895
      ("1001001101010001", '0', '1', "01", "101", "001", "011", '0', '-', "00"), -- i=4896
      ("1001101101010001", '1', '1', "01", "101", "001", "011", '0', '-', "00"), -- i=4897
      ("1001101101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4898
      ("1010001101010001", '0', '1', "10", "101", "001", "011", '0', '-', "00"), -- i=4899
      ("1010101101010001", '1', '1', "10", "101", "001", "011", '0', '-', "00"), -- i=4900
      ("1010101101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4901
      ("1011001101010001", '0', '1', "11", "101", "001", "011", '0', '-', "00"), -- i=4902
      ("1011101101010001", '1', '1', "11", "101", "001", "011", '0', '-', "00"), -- i=4903
      ("1011101101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4904
      ("0101001101010000", '0', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=4905
      ("0101101101010000", '1', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=4906
      ("0101101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4907
      ("0100001101010000", '0', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=4908
      ("0100101101010000", '1', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=4909
      ("0100101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4910
      ("0000001111100100", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4911
      ("0000101111100100", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4912
      ("0000101111100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4913
      ("1000001101010010", '0', '1', "00", "101", "010", "011", '0', '-', "00"), -- i=4914
      ("1000101101010010", '1', '1', "00", "101", "010", "011", '0', '-', "00"), -- i=4915
      ("1000101101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4916
      ("1001001101010010", '0', '1', "01", "101", "010", "011", '0', '-', "00"), -- i=4917
      ("1001101101010010", '1', '1', "01", "101", "010", "011", '0', '-', "00"), -- i=4918
      ("1001101101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4919
      ("1010001101010010", '0', '1', "10", "101", "010", "011", '0', '-', "00"), -- i=4920
      ("1010101101010010", '1', '1', "10", "101", "010", "011", '0', '-', "00"), -- i=4921
      ("1010101101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4922
      ("1011001101010010", '0', '1', "11", "101", "010", "011", '0', '-', "00"), -- i=4923
      ("1011101101010010", '1', '1', "11", "101", "010", "011", '0', '-', "00"), -- i=4924
      ("1011101101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4925
      ("0101001101010000", '0', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=4926
      ("0101101101010000", '1', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=4927
      ("0101101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4928
      ("0100001101010000", '0', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=4929
      ("0100101101010000", '1', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=4930
      ("0100101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4931
      ("0000001100010010", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4932
      ("0000101100010010", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4933
      ("0000101100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4934
      ("1000001101010011", '0', '1', "00", "101", "011", "011", '0', '-', "00"), -- i=4935
      ("1000101101010011", '1', '1', "00", "101", "011", "011", '0', '-', "00"), -- i=4936
      ("1000101101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4937
      ("1001001101010011", '0', '1', "01", "101", "011", "011", '0', '-', "00"), -- i=4938
      ("1001101101010011", '1', '1', "01", "101", "011", "011", '0', '-', "00"), -- i=4939
      ("1001101101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4940
      ("1010001101010011", '0', '1', "10", "101", "011", "011", '0', '-', "00"), -- i=4941
      ("1010101101010011", '1', '1', "10", "101", "011", "011", '0', '-', "00"), -- i=4942
      ("1010101101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4943
      ("1011001101010011", '0', '1', "11", "101", "011", "011", '0', '-', "00"), -- i=4944
      ("1011101101010011", '1', '1', "11", "101", "011", "011", '0', '-', "00"), -- i=4945
      ("1011101101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4946
      ("0101001101010000", '0', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=4947
      ("0101101101010000", '1', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=4948
      ("0101101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4949
      ("0100001101010000", '0', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=4950
      ("0100101101010000", '1', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=4951
      ("0100101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4952
      ("0000001110000001", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4953
      ("0000101110000001", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4954
      ("0000101110000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4955
      ("1000001101010100", '0', '1', "00", "101", "100", "011", '0', '-', "00"), -- i=4956
      ("1000101101010100", '1', '1', "00", "101", "100", "011", '0', '-', "00"), -- i=4957
      ("1000101101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4958
      ("1001001101010100", '0', '1', "01", "101", "100", "011", '0', '-', "00"), -- i=4959
      ("1001101101010100", '1', '1', "01", "101", "100", "011", '0', '-', "00"), -- i=4960
      ("1001101101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4961
      ("1010001101010100", '0', '1', "10", "101", "100", "011", '0', '-', "00"), -- i=4962
      ("1010101101010100", '1', '1', "10", "101", "100", "011", '0', '-', "00"), -- i=4963
      ("1010101101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4964
      ("1011001101010100", '0', '1', "11", "101", "100", "011", '0', '-', "00"), -- i=4965
      ("1011101101010100", '1', '1', "11", "101", "100", "011", '0', '-', "00"), -- i=4966
      ("1011101101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4967
      ("0101001101010000", '0', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=4968
      ("0101101101010000", '1', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=4969
      ("0101101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4970
      ("0100001101010000", '0', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=4971
      ("0100101101010000", '1', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=4972
      ("0100101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4973
      ("0000001111000010", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4974
      ("0000101111000010", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4975
      ("0000101111000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4976
      ("1000001101010101", '0', '1', "00", "101", "101", "011", '0', '-', "00"), -- i=4977
      ("1000101101010101", '1', '1', "00", "101", "101", "011", '0', '-', "00"), -- i=4978
      ("1000101101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4979
      ("1001001101010101", '0', '1', "01", "101", "101", "011", '0', '-', "00"), -- i=4980
      ("1001101101010101", '1', '1', "01", "101", "101", "011", '0', '-', "00"), -- i=4981
      ("1001101101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4982
      ("1010001101010101", '0', '1', "10", "101", "101", "011", '0', '-', "00"), -- i=4983
      ("1010101101010101", '1', '1', "10", "101", "101", "011", '0', '-', "00"), -- i=4984
      ("1010101101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4985
      ("1011001101010101", '0', '1', "11", "101", "101", "011", '0', '-', "00"), -- i=4986
      ("1011101101010101", '1', '1', "11", "101", "101", "011", '0', '-', "00"), -- i=4987
      ("1011101101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4988
      ("0101001101010000", '0', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=4989
      ("0101101101010000", '1', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=4990
      ("0101101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4991
      ("0100001101010000", '0', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=4992
      ("0100101101010000", '1', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=4993
      ("0100101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4994
      ("0000001111010000", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4995
      ("0000101111010000", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=4996
      ("0000101111010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=4997
      ("1000001101010110", '0', '1', "00", "101", "110", "011", '0', '-', "00"), -- i=4998
      ("1000101101010110", '1', '1', "00", "101", "110", "011", '0', '-', "00"), -- i=4999
      ("1000101101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5000
      ("1001001101010110", '0', '1', "01", "101", "110", "011", '0', '-', "00"), -- i=5001
      ("1001101101010110", '1', '1', "01", "101", "110", "011", '0', '-', "00"), -- i=5002
      ("1001101101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5003
      ("1010001101010110", '0', '1', "10", "101", "110", "011", '0', '-', "00"), -- i=5004
      ("1010101101010110", '1', '1', "10", "101", "110", "011", '0', '-', "00"), -- i=5005
      ("1010101101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5006
      ("1011001101010110", '0', '1', "11", "101", "110", "011", '0', '-', "00"), -- i=5007
      ("1011101101010110", '1', '1', "11", "101", "110", "011", '0', '-', "00"), -- i=5008
      ("1011101101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5009
      ("0101001101010000", '0', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=5010
      ("0101101101010000", '1', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=5011
      ("0101101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5012
      ("0100001101010000", '0', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=5013
      ("0100101101010000", '1', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=5014
      ("0100101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5015
      ("0000001100001011", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5016
      ("0000101100001011", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5017
      ("0000101100001011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5018
      ("1000001101010111", '0', '1', "00", "101", "111", "011", '0', '-', "00"), -- i=5019
      ("1000101101010111", '1', '1', "00", "101", "111", "011", '0', '-', "00"), -- i=5020
      ("1000101101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5021
      ("1001001101010111", '0', '1', "01", "101", "111", "011", '0', '-', "00"), -- i=5022
      ("1001101101010111", '1', '1', "01", "101", "111", "011", '0', '-', "00"), -- i=5023
      ("1001101101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5024
      ("1010001101010111", '0', '1', "10", "101", "111", "011", '0', '-', "00"), -- i=5025
      ("1010101101010111", '1', '1', "10", "101", "111", "011", '0', '-', "00"), -- i=5026
      ("1010101101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5027
      ("1011001101010111", '0', '1', "11", "101", "111", "011", '0', '-', "00"), -- i=5028
      ("1011101101010111", '1', '1', "11", "101", "111", "011", '0', '-', "00"), -- i=5029
      ("1011101101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5030
      ("0101001101010000", '0', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=5031
      ("0101101101010000", '1', '1', "--", "101", "---", "011", '0', '1', "01"), -- i=5032
      ("0101101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5033
      ("0100001101010000", '0', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=5034
      ("0100101101010000", '1', '0', "--", "101", "011", "---", '1', '-', "--"), -- i=5035
      ("0100101101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5036
      ("0000001100000101", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5037
      ("0000101100000101", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5038
      ("0000101100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5039
      ("1000001101100000", '0', '1', "00", "110", "000", "011", '0', '-', "00"), -- i=5040
      ("1000101101100000", '1', '1', "00", "110", "000", "011", '0', '-', "00"), -- i=5041
      ("1000101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5042
      ("1001001101100000", '0', '1', "01", "110", "000", "011", '0', '-', "00"), -- i=5043
      ("1001101101100000", '1', '1', "01", "110", "000", "011", '0', '-', "00"), -- i=5044
      ("1001101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5045
      ("1010001101100000", '0', '1', "10", "110", "000", "011", '0', '-', "00"), -- i=5046
      ("1010101101100000", '1', '1', "10", "110", "000", "011", '0', '-', "00"), -- i=5047
      ("1010101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5048
      ("1011001101100000", '0', '1', "11", "110", "000", "011", '0', '-', "00"), -- i=5049
      ("1011101101100000", '1', '1', "11", "110", "000", "011", '0', '-', "00"), -- i=5050
      ("1011101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5051
      ("0101001101100000", '0', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5052
      ("0101101101100000", '1', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5053
      ("0101101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5054
      ("0100001101100000", '0', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5055
      ("0100101101100000", '1', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5056
      ("0100101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5057
      ("0000001100011011", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5058
      ("0000101100011011", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5059
      ("0000101100011011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5060
      ("1000001101100001", '0', '1', "00", "110", "001", "011", '0', '-', "00"), -- i=5061
      ("1000101101100001", '1', '1', "00", "110", "001", "011", '0', '-', "00"), -- i=5062
      ("1000101101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5063
      ("1001001101100001", '0', '1', "01", "110", "001", "011", '0', '-', "00"), -- i=5064
      ("1001101101100001", '1', '1', "01", "110", "001", "011", '0', '-', "00"), -- i=5065
      ("1001101101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5066
      ("1010001101100001", '0', '1', "10", "110", "001", "011", '0', '-', "00"), -- i=5067
      ("1010101101100001", '1', '1', "10", "110", "001", "011", '0', '-', "00"), -- i=5068
      ("1010101101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5069
      ("1011001101100001", '0', '1', "11", "110", "001", "011", '0', '-', "00"), -- i=5070
      ("1011101101100001", '1', '1', "11", "110", "001", "011", '0', '-', "00"), -- i=5071
      ("1011101101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5072
      ("0101001101100000", '0', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5073
      ("0101101101100000", '1', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5074
      ("0101101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5075
      ("0100001101100000", '0', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5076
      ("0100101101100000", '1', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5077
      ("0100101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5078
      ("0000001110000010", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5079
      ("0000101110000010", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5080
      ("0000101110000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5081
      ("1000001101100010", '0', '1', "00", "110", "010", "011", '0', '-', "00"), -- i=5082
      ("1000101101100010", '1', '1', "00", "110", "010", "011", '0', '-', "00"), -- i=5083
      ("1000101101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5084
      ("1001001101100010", '0', '1', "01", "110", "010", "011", '0', '-', "00"), -- i=5085
      ("1001101101100010", '1', '1', "01", "110", "010", "011", '0', '-', "00"), -- i=5086
      ("1001101101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5087
      ("1010001101100010", '0', '1', "10", "110", "010", "011", '0', '-', "00"), -- i=5088
      ("1010101101100010", '1', '1', "10", "110", "010", "011", '0', '-', "00"), -- i=5089
      ("1010101101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5090
      ("1011001101100010", '0', '1', "11", "110", "010", "011", '0', '-', "00"), -- i=5091
      ("1011101101100010", '1', '1', "11", "110", "010", "011", '0', '-', "00"), -- i=5092
      ("1011101101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5093
      ("0101001101100000", '0', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5094
      ("0101101101100000", '1', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5095
      ("0101101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5096
      ("0100001101100000", '0', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5097
      ("0100101101100000", '1', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5098
      ("0100101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5099
      ("0000001110010110", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5100
      ("0000101110010110", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5101
      ("0000101110010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5102
      ("1000001101100011", '0', '1', "00", "110", "011", "011", '0', '-', "00"), -- i=5103
      ("1000101101100011", '1', '1', "00", "110", "011", "011", '0', '-', "00"), -- i=5104
      ("1000101101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5105
      ("1001001101100011", '0', '1', "01", "110", "011", "011", '0', '-', "00"), -- i=5106
      ("1001101101100011", '1', '1', "01", "110", "011", "011", '0', '-', "00"), -- i=5107
      ("1001101101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5108
      ("1010001101100011", '0', '1', "10", "110", "011", "011", '0', '-', "00"), -- i=5109
      ("1010101101100011", '1', '1', "10", "110", "011", "011", '0', '-', "00"), -- i=5110
      ("1010101101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5111
      ("1011001101100011", '0', '1', "11", "110", "011", "011", '0', '-', "00"), -- i=5112
      ("1011101101100011", '1', '1', "11", "110", "011", "011", '0', '-', "00"), -- i=5113
      ("1011101101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5114
      ("0101001101100000", '0', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5115
      ("0101101101100000", '1', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5116
      ("0101101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5117
      ("0100001101100000", '0', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5118
      ("0100101101100000", '1', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5119
      ("0100101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5120
      ("0000001101001111", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5121
      ("0000101101001111", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5122
      ("0000101101001111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5123
      ("1000001101100100", '0', '1', "00", "110", "100", "011", '0', '-', "00"), -- i=5124
      ("1000101101100100", '1', '1', "00", "110", "100", "011", '0', '-', "00"), -- i=5125
      ("1000101101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5126
      ("1001001101100100", '0', '1', "01", "110", "100", "011", '0', '-', "00"), -- i=5127
      ("1001101101100100", '1', '1', "01", "110", "100", "011", '0', '-', "00"), -- i=5128
      ("1001101101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5129
      ("1010001101100100", '0', '1', "10", "110", "100", "011", '0', '-', "00"), -- i=5130
      ("1010101101100100", '1', '1', "10", "110", "100", "011", '0', '-', "00"), -- i=5131
      ("1010101101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5132
      ("1011001101100100", '0', '1', "11", "110", "100", "011", '0', '-', "00"), -- i=5133
      ("1011101101100100", '1', '1', "11", "110", "100", "011", '0', '-', "00"), -- i=5134
      ("1011101101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5135
      ("0101001101100000", '0', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5136
      ("0101101101100000", '1', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5137
      ("0101101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5138
      ("0100001101100000", '0', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5139
      ("0100101101100000", '1', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5140
      ("0100101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5141
      ("0000001111110111", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5142
      ("0000101111110111", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5143
      ("0000101111110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5144
      ("1000001101100101", '0', '1', "00", "110", "101", "011", '0', '-', "00"), -- i=5145
      ("1000101101100101", '1', '1', "00", "110", "101", "011", '0', '-', "00"), -- i=5146
      ("1000101101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5147
      ("1001001101100101", '0', '1', "01", "110", "101", "011", '0', '-', "00"), -- i=5148
      ("1001101101100101", '1', '1', "01", "110", "101", "011", '0', '-', "00"), -- i=5149
      ("1001101101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5150
      ("1010001101100101", '0', '1', "10", "110", "101", "011", '0', '-', "00"), -- i=5151
      ("1010101101100101", '1', '1', "10", "110", "101", "011", '0', '-', "00"), -- i=5152
      ("1010101101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5153
      ("1011001101100101", '0', '1', "11", "110", "101", "011", '0', '-', "00"), -- i=5154
      ("1011101101100101", '1', '1', "11", "110", "101", "011", '0', '-', "00"), -- i=5155
      ("1011101101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5156
      ("0101001101100000", '0', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5157
      ("0101101101100000", '1', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5158
      ("0101101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5159
      ("0100001101100000", '0', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5160
      ("0100101101100000", '1', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5161
      ("0100101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5162
      ("0000001101000010", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5163
      ("0000101101000010", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5164
      ("0000101101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5165
      ("1000001101100110", '0', '1', "00", "110", "110", "011", '0', '-', "00"), -- i=5166
      ("1000101101100110", '1', '1', "00", "110", "110", "011", '0', '-', "00"), -- i=5167
      ("1000101101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5168
      ("1001001101100110", '0', '1', "01", "110", "110", "011", '0', '-', "00"), -- i=5169
      ("1001101101100110", '1', '1', "01", "110", "110", "011", '0', '-', "00"), -- i=5170
      ("1001101101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5171
      ("1010001101100110", '0', '1', "10", "110", "110", "011", '0', '-', "00"), -- i=5172
      ("1010101101100110", '1', '1', "10", "110", "110", "011", '0', '-', "00"), -- i=5173
      ("1010101101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5174
      ("1011001101100110", '0', '1', "11", "110", "110", "011", '0', '-', "00"), -- i=5175
      ("1011101101100110", '1', '1', "11", "110", "110", "011", '0', '-', "00"), -- i=5176
      ("1011101101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5177
      ("0101001101100000", '0', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5178
      ("0101101101100000", '1', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5179
      ("0101101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5180
      ("0100001101100000", '0', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5181
      ("0100101101100000", '1', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5182
      ("0100101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5183
      ("0000001111001111", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5184
      ("0000101111001111", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5185
      ("0000101111001111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5186
      ("1000001101100111", '0', '1', "00", "110", "111", "011", '0', '-', "00"), -- i=5187
      ("1000101101100111", '1', '1', "00", "110", "111", "011", '0', '-', "00"), -- i=5188
      ("1000101101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5189
      ("1001001101100111", '0', '1', "01", "110", "111", "011", '0', '-', "00"), -- i=5190
      ("1001101101100111", '1', '1', "01", "110", "111", "011", '0', '-', "00"), -- i=5191
      ("1001101101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5192
      ("1010001101100111", '0', '1', "10", "110", "111", "011", '0', '-', "00"), -- i=5193
      ("1010101101100111", '1', '1', "10", "110", "111", "011", '0', '-', "00"), -- i=5194
      ("1010101101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5195
      ("1011001101100111", '0', '1', "11", "110", "111", "011", '0', '-', "00"), -- i=5196
      ("1011101101100111", '1', '1', "11", "110", "111", "011", '0', '-', "00"), -- i=5197
      ("1011101101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5198
      ("0101001101100000", '0', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5199
      ("0101101101100000", '1', '1', "--", "110", "---", "011", '0', '1', "01"), -- i=5200
      ("0101101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5201
      ("0100001101100000", '0', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5202
      ("0100101101100000", '1', '0', "--", "110", "011", "---", '1', '-', "--"), -- i=5203
      ("0100101101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5204
      ("0000001110001111", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5205
      ("0000101110001111", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5206
      ("0000101110001111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5207
      ("1000001101110000", '0', '1', "00", "111", "000", "011", '0', '-', "00"), -- i=5208
      ("1000101101110000", '1', '1', "00", "111", "000", "011", '0', '-', "00"), -- i=5209
      ("1000101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5210
      ("1001001101110000", '0', '1', "01", "111", "000", "011", '0', '-', "00"), -- i=5211
      ("1001101101110000", '1', '1', "01", "111", "000", "011", '0', '-', "00"), -- i=5212
      ("1001101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5213
      ("1010001101110000", '0', '1', "10", "111", "000", "011", '0', '-', "00"), -- i=5214
      ("1010101101110000", '1', '1', "10", "111", "000", "011", '0', '-', "00"), -- i=5215
      ("1010101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5216
      ("1011001101110000", '0', '1', "11", "111", "000", "011", '0', '-', "00"), -- i=5217
      ("1011101101110000", '1', '1', "11", "111", "000", "011", '0', '-', "00"), -- i=5218
      ("1011101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5219
      ("0101001101110000", '0', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5220
      ("0101101101110000", '1', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5221
      ("0101101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5222
      ("0100001101110000", '0', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5223
      ("0100101101110000", '1', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5224
      ("0100101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5225
      ("0000001101111111", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5226
      ("0000101101111111", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5227
      ("0000101101111111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5228
      ("1000001101110001", '0', '1', "00", "111", "001", "011", '0', '-', "00"), -- i=5229
      ("1000101101110001", '1', '1', "00", "111", "001", "011", '0', '-', "00"), -- i=5230
      ("1000101101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5231
      ("1001001101110001", '0', '1', "01", "111", "001", "011", '0', '-', "00"), -- i=5232
      ("1001101101110001", '1', '1', "01", "111", "001", "011", '0', '-', "00"), -- i=5233
      ("1001101101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5234
      ("1010001101110001", '0', '1', "10", "111", "001", "011", '0', '-', "00"), -- i=5235
      ("1010101101110001", '1', '1', "10", "111", "001", "011", '0', '-', "00"), -- i=5236
      ("1010101101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5237
      ("1011001101110001", '0', '1', "11", "111", "001", "011", '0', '-', "00"), -- i=5238
      ("1011101101110001", '1', '1', "11", "111", "001", "011", '0', '-', "00"), -- i=5239
      ("1011101101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5240
      ("0101001101110000", '0', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5241
      ("0101101101110000", '1', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5242
      ("0101101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5243
      ("0100001101110000", '0', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5244
      ("0100101101110000", '1', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5245
      ("0100101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5246
      ("0000001111001110", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5247
      ("0000101111001110", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5248
      ("0000101111001110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5249
      ("1000001101110010", '0', '1', "00", "111", "010", "011", '0', '-', "00"), -- i=5250
      ("1000101101110010", '1', '1', "00", "111", "010", "011", '0', '-', "00"), -- i=5251
      ("1000101101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5252
      ("1001001101110010", '0', '1', "01", "111", "010", "011", '0', '-', "00"), -- i=5253
      ("1001101101110010", '1', '1', "01", "111", "010", "011", '0', '-', "00"), -- i=5254
      ("1001101101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5255
      ("1010001101110010", '0', '1', "10", "111", "010", "011", '0', '-', "00"), -- i=5256
      ("1010101101110010", '1', '1', "10", "111", "010", "011", '0', '-', "00"), -- i=5257
      ("1010101101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5258
      ("1011001101110010", '0', '1', "11", "111", "010", "011", '0', '-', "00"), -- i=5259
      ("1011101101110010", '1', '1', "11", "111", "010", "011", '0', '-', "00"), -- i=5260
      ("1011101101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5261
      ("0101001101110000", '0', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5262
      ("0101101101110000", '1', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5263
      ("0101101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5264
      ("0100001101110000", '0', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5265
      ("0100101101110000", '1', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5266
      ("0100101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5267
      ("0000001101010111", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5268
      ("0000101101010111", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5269
      ("0000101101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5270
      ("1000001101110011", '0', '1', "00", "111", "011", "011", '0', '-', "00"), -- i=5271
      ("1000101101110011", '1', '1', "00", "111", "011", "011", '0', '-', "00"), -- i=5272
      ("1000101101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5273
      ("1001001101110011", '0', '1', "01", "111", "011", "011", '0', '-', "00"), -- i=5274
      ("1001101101110011", '1', '1', "01", "111", "011", "011", '0', '-', "00"), -- i=5275
      ("1001101101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5276
      ("1010001101110011", '0', '1', "10", "111", "011", "011", '0', '-', "00"), -- i=5277
      ("1010101101110011", '1', '1', "10", "111", "011", "011", '0', '-', "00"), -- i=5278
      ("1010101101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5279
      ("1011001101110011", '0', '1', "11", "111", "011", "011", '0', '-', "00"), -- i=5280
      ("1011101101110011", '1', '1', "11", "111", "011", "011", '0', '-', "00"), -- i=5281
      ("1011101101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5282
      ("0101001101110000", '0', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5283
      ("0101101101110000", '1', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5284
      ("0101101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5285
      ("0100001101110000", '0', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5286
      ("0100101101110000", '1', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5287
      ("0100101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5288
      ("0000001110000100", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5289
      ("0000101110000100", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5290
      ("0000101110000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5291
      ("1000001101110100", '0', '1', "00", "111", "100", "011", '0', '-', "00"), -- i=5292
      ("1000101101110100", '1', '1', "00", "111", "100", "011", '0', '-', "00"), -- i=5293
      ("1000101101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5294
      ("1001001101110100", '0', '1', "01", "111", "100", "011", '0', '-', "00"), -- i=5295
      ("1001101101110100", '1', '1', "01", "111", "100", "011", '0', '-', "00"), -- i=5296
      ("1001101101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5297
      ("1010001101110100", '0', '1', "10", "111", "100", "011", '0', '-', "00"), -- i=5298
      ("1010101101110100", '1', '1', "10", "111", "100", "011", '0', '-', "00"), -- i=5299
      ("1010101101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5300
      ("1011001101110100", '0', '1', "11", "111", "100", "011", '0', '-', "00"), -- i=5301
      ("1011101101110100", '1', '1', "11", "111", "100", "011", '0', '-', "00"), -- i=5302
      ("1011101101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5303
      ("0101001101110000", '0', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5304
      ("0101101101110000", '1', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5305
      ("0101101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5306
      ("0100001101110000", '0', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5307
      ("0100101101110000", '1', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5308
      ("0100101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5309
      ("0000001100100110", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5310
      ("0000101100100110", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5311
      ("0000101100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5312
      ("1000001101110101", '0', '1', "00", "111", "101", "011", '0', '-', "00"), -- i=5313
      ("1000101101110101", '1', '1', "00", "111", "101", "011", '0', '-', "00"), -- i=5314
      ("1000101101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5315
      ("1001001101110101", '0', '1', "01", "111", "101", "011", '0', '-', "00"), -- i=5316
      ("1001101101110101", '1', '1', "01", "111", "101", "011", '0', '-', "00"), -- i=5317
      ("1001101101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5318
      ("1010001101110101", '0', '1', "10", "111", "101", "011", '0', '-', "00"), -- i=5319
      ("1010101101110101", '1', '1', "10", "111", "101", "011", '0', '-', "00"), -- i=5320
      ("1010101101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5321
      ("1011001101110101", '0', '1', "11", "111", "101", "011", '0', '-', "00"), -- i=5322
      ("1011101101110101", '1', '1', "11", "111", "101", "011", '0', '-', "00"), -- i=5323
      ("1011101101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5324
      ("0101001101110000", '0', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5325
      ("0101101101110000", '1', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5326
      ("0101101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5327
      ("0100001101110000", '0', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5328
      ("0100101101110000", '1', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5329
      ("0100101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5330
      ("0000001101111101", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5331
      ("0000101101111101", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5332
      ("0000101101111101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5333
      ("1000001101110110", '0', '1', "00", "111", "110", "011", '0', '-', "00"), -- i=5334
      ("1000101101110110", '1', '1', "00", "111", "110", "011", '0', '-', "00"), -- i=5335
      ("1000101101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5336
      ("1001001101110110", '0', '1', "01", "111", "110", "011", '0', '-', "00"), -- i=5337
      ("1001101101110110", '1', '1', "01", "111", "110", "011", '0', '-', "00"), -- i=5338
      ("1001101101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5339
      ("1010001101110110", '0', '1', "10", "111", "110", "011", '0', '-', "00"), -- i=5340
      ("1010101101110110", '1', '1', "10", "111", "110", "011", '0', '-', "00"), -- i=5341
      ("1010101101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5342
      ("1011001101110110", '0', '1', "11", "111", "110", "011", '0', '-', "00"), -- i=5343
      ("1011101101110110", '1', '1', "11", "111", "110", "011", '0', '-', "00"), -- i=5344
      ("1011101101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5345
      ("0101001101110000", '0', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5346
      ("0101101101110000", '1', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5347
      ("0101101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5348
      ("0100001101110000", '0', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5349
      ("0100101101110000", '1', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5350
      ("0100101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5351
      ("0000001100011101", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5352
      ("0000101100011101", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5353
      ("0000101100011101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5354
      ("1000001101110111", '0', '1', "00", "111", "111", "011", '0', '-', "00"), -- i=5355
      ("1000101101110111", '1', '1', "00", "111", "111", "011", '0', '-', "00"), -- i=5356
      ("1000101101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5357
      ("1001001101110111", '0', '1', "01", "111", "111", "011", '0', '-', "00"), -- i=5358
      ("1001101101110111", '1', '1', "01", "111", "111", "011", '0', '-', "00"), -- i=5359
      ("1001101101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5360
      ("1010001101110111", '0', '1', "10", "111", "111", "011", '0', '-', "00"), -- i=5361
      ("1010101101110111", '1', '1', "10", "111", "111", "011", '0', '-', "00"), -- i=5362
      ("1010101101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5363
      ("1011001101110111", '0', '1', "11", "111", "111", "011", '0', '-', "00"), -- i=5364
      ("1011101101110111", '1', '1', "11", "111", "111", "011", '0', '-', "00"), -- i=5365
      ("1011101101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5366
      ("0101001101110000", '0', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5367
      ("0101101101110000", '1', '1', "--", "111", "---", "011", '0', '1', "01"), -- i=5368
      ("0101101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5369
      ("0100001101110000", '0', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5370
      ("0100101101110000", '1', '0', "--", "111", "011", "---", '1', '-', "--"), -- i=5371
      ("0100101101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5372
      ("0000001101010110", '0', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5373
      ("0000101101010110", '1', '1', "--", "---", "---", "011", '0', '-', "10"), -- i=5374
      ("0000101101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5375
      ("1000010000000000", '0', '1', "00", "000", "000", "100", '0', '-', "00"), -- i=5376
      ("1000110000000000", '1', '1', "00", "000", "000", "100", '0', '-', "00"), -- i=5377
      ("1000110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5378
      ("1001010000000000", '0', '1', "01", "000", "000", "100", '0', '-', "00"), -- i=5379
      ("1001110000000000", '1', '1', "01", "000", "000", "100", '0', '-', "00"), -- i=5380
      ("1001110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5381
      ("1010010000000000", '0', '1', "10", "000", "000", "100", '0', '-', "00"), -- i=5382
      ("1010110000000000", '1', '1', "10", "000", "000", "100", '0', '-', "00"), -- i=5383
      ("1010110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5384
      ("1011010000000000", '0', '1', "11", "000", "000", "100", '0', '-', "00"), -- i=5385
      ("1011110000000000", '1', '1', "11", "000", "000", "100", '0', '-', "00"), -- i=5386
      ("1011110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5387
      ("0101010000000000", '0', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5388
      ("0101110000000000", '1', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5389
      ("0101110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5390
      ("0100010000000000", '0', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5391
      ("0100110000000000", '1', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5392
      ("0100110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5393
      ("0000010000000111", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5394
      ("0000110000000111", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5395
      ("0000110000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5396
      ("1000010000000001", '0', '1', "00", "000", "001", "100", '0', '-', "00"), -- i=5397
      ("1000110000000001", '1', '1', "00", "000", "001", "100", '0', '-', "00"), -- i=5398
      ("1000110000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5399
      ("1001010000000001", '0', '1', "01", "000", "001", "100", '0', '-', "00"), -- i=5400
      ("1001110000000001", '1', '1', "01", "000", "001", "100", '0', '-', "00"), -- i=5401
      ("1001110000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5402
      ("1010010000000001", '0', '1', "10", "000", "001", "100", '0', '-', "00"), -- i=5403
      ("1010110000000001", '1', '1', "10", "000", "001", "100", '0', '-', "00"), -- i=5404
      ("1010110000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5405
      ("1011010000000001", '0', '1', "11", "000", "001", "100", '0', '-', "00"), -- i=5406
      ("1011110000000001", '1', '1', "11", "000", "001", "100", '0', '-', "00"), -- i=5407
      ("1011110000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5408
      ("0101010000000000", '0', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5409
      ("0101110000000000", '1', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5410
      ("0101110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5411
      ("0100010000000000", '0', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5412
      ("0100110000000000", '1', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5413
      ("0100110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5414
      ("0000010000101100", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5415
      ("0000110000101100", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5416
      ("0000110000101100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5417
      ("1000010000000010", '0', '1', "00", "000", "010", "100", '0', '-', "00"), -- i=5418
      ("1000110000000010", '1', '1', "00", "000", "010", "100", '0', '-', "00"), -- i=5419
      ("1000110000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5420
      ("1001010000000010", '0', '1', "01", "000", "010", "100", '0', '-', "00"), -- i=5421
      ("1001110000000010", '1', '1', "01", "000", "010", "100", '0', '-', "00"), -- i=5422
      ("1001110000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5423
      ("1010010000000010", '0', '1', "10", "000", "010", "100", '0', '-', "00"), -- i=5424
      ("1010110000000010", '1', '1', "10", "000", "010", "100", '0', '-', "00"), -- i=5425
      ("1010110000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5426
      ("1011010000000010", '0', '1', "11", "000", "010", "100", '0', '-', "00"), -- i=5427
      ("1011110000000010", '1', '1', "11", "000", "010", "100", '0', '-', "00"), -- i=5428
      ("1011110000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5429
      ("0101010000000000", '0', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5430
      ("0101110000000000", '1', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5431
      ("0101110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5432
      ("0100010000000000", '0', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5433
      ("0100110000000000", '1', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5434
      ("0100110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5435
      ("0000010000101000", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5436
      ("0000110000101000", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5437
      ("0000110000101000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5438
      ("1000010000000011", '0', '1', "00", "000", "011", "100", '0', '-', "00"), -- i=5439
      ("1000110000000011", '1', '1', "00", "000", "011", "100", '0', '-', "00"), -- i=5440
      ("1000110000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5441
      ("1001010000000011", '0', '1', "01", "000", "011", "100", '0', '-', "00"), -- i=5442
      ("1001110000000011", '1', '1', "01", "000", "011", "100", '0', '-', "00"), -- i=5443
      ("1001110000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5444
      ("1010010000000011", '0', '1', "10", "000", "011", "100", '0', '-', "00"), -- i=5445
      ("1010110000000011", '1', '1', "10", "000", "011", "100", '0', '-', "00"), -- i=5446
      ("1010110000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5447
      ("1011010000000011", '0', '1', "11", "000", "011", "100", '0', '-', "00"), -- i=5448
      ("1011110000000011", '1', '1', "11", "000", "011", "100", '0', '-', "00"), -- i=5449
      ("1011110000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5450
      ("0101010000000000", '0', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5451
      ("0101110000000000", '1', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5452
      ("0101110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5453
      ("0100010000000000", '0', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5454
      ("0100110000000000", '1', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5455
      ("0100110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5456
      ("0000010001111110", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5457
      ("0000110001111110", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5458
      ("0000110001111110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5459
      ("1000010000000100", '0', '1', "00", "000", "100", "100", '0', '-', "00"), -- i=5460
      ("1000110000000100", '1', '1', "00", "000", "100", "100", '0', '-', "00"), -- i=5461
      ("1000110000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5462
      ("1001010000000100", '0', '1', "01", "000", "100", "100", '0', '-', "00"), -- i=5463
      ("1001110000000100", '1', '1', "01", "000", "100", "100", '0', '-', "00"), -- i=5464
      ("1001110000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5465
      ("1010010000000100", '0', '1', "10", "000", "100", "100", '0', '-', "00"), -- i=5466
      ("1010110000000100", '1', '1', "10", "000", "100", "100", '0', '-', "00"), -- i=5467
      ("1010110000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5468
      ("1011010000000100", '0', '1', "11", "000", "100", "100", '0', '-', "00"), -- i=5469
      ("1011110000000100", '1', '1', "11", "000", "100", "100", '0', '-', "00"), -- i=5470
      ("1011110000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5471
      ("0101010000000000", '0', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5472
      ("0101110000000000", '1', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5473
      ("0101110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5474
      ("0100010000000000", '0', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5475
      ("0100110000000000", '1', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5476
      ("0100110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5477
      ("0000010001011111", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5478
      ("0000110001011111", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5479
      ("0000110001011111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5480
      ("1000010000000101", '0', '1', "00", "000", "101", "100", '0', '-', "00"), -- i=5481
      ("1000110000000101", '1', '1', "00", "000", "101", "100", '0', '-', "00"), -- i=5482
      ("1000110000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5483
      ("1001010000000101", '0', '1', "01", "000", "101", "100", '0', '-', "00"), -- i=5484
      ("1001110000000101", '1', '1', "01", "000", "101", "100", '0', '-', "00"), -- i=5485
      ("1001110000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5486
      ("1010010000000101", '0', '1', "10", "000", "101", "100", '0', '-', "00"), -- i=5487
      ("1010110000000101", '1', '1', "10", "000", "101", "100", '0', '-', "00"), -- i=5488
      ("1010110000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5489
      ("1011010000000101", '0', '1', "11", "000", "101", "100", '0', '-', "00"), -- i=5490
      ("1011110000000101", '1', '1', "11", "000", "101", "100", '0', '-', "00"), -- i=5491
      ("1011110000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5492
      ("0101010000000000", '0', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5493
      ("0101110000000000", '1', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5494
      ("0101110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5495
      ("0100010000000000", '0', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5496
      ("0100110000000000", '1', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5497
      ("0100110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5498
      ("0000010011011111", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5499
      ("0000110011011111", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5500
      ("0000110011011111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5501
      ("1000010000000110", '0', '1', "00", "000", "110", "100", '0', '-', "00"), -- i=5502
      ("1000110000000110", '1', '1', "00", "000", "110", "100", '0', '-', "00"), -- i=5503
      ("1000110000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5504
      ("1001010000000110", '0', '1', "01", "000", "110", "100", '0', '-', "00"), -- i=5505
      ("1001110000000110", '1', '1', "01", "000", "110", "100", '0', '-', "00"), -- i=5506
      ("1001110000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5507
      ("1010010000000110", '0', '1', "10", "000", "110", "100", '0', '-', "00"), -- i=5508
      ("1010110000000110", '1', '1', "10", "000", "110", "100", '0', '-', "00"), -- i=5509
      ("1010110000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5510
      ("1011010000000110", '0', '1', "11", "000", "110", "100", '0', '-', "00"), -- i=5511
      ("1011110000000110", '1', '1', "11", "000", "110", "100", '0', '-', "00"), -- i=5512
      ("1011110000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5513
      ("0101010000000000", '0', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5514
      ("0101110000000000", '1', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5515
      ("0101110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5516
      ("0100010000000000", '0', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5517
      ("0100110000000000", '1', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5518
      ("0100110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5519
      ("0000010000110001", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5520
      ("0000110000110001", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5521
      ("0000110000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5522
      ("1000010000000111", '0', '1', "00", "000", "111", "100", '0', '-', "00"), -- i=5523
      ("1000110000000111", '1', '1', "00", "000", "111", "100", '0', '-', "00"), -- i=5524
      ("1000110000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5525
      ("1001010000000111", '0', '1', "01", "000", "111", "100", '0', '-', "00"), -- i=5526
      ("1001110000000111", '1', '1', "01", "000", "111", "100", '0', '-', "00"), -- i=5527
      ("1001110000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5528
      ("1010010000000111", '0', '1', "10", "000", "111", "100", '0', '-', "00"), -- i=5529
      ("1010110000000111", '1', '1', "10", "000", "111", "100", '0', '-', "00"), -- i=5530
      ("1010110000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5531
      ("1011010000000111", '0', '1', "11", "000", "111", "100", '0', '-', "00"), -- i=5532
      ("1011110000000111", '1', '1', "11", "000", "111", "100", '0', '-', "00"), -- i=5533
      ("1011110000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5534
      ("0101010000000000", '0', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5535
      ("0101110000000000", '1', '1', "--", "000", "---", "100", '0', '1', "01"), -- i=5536
      ("0101110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5537
      ("0100010000000000", '0', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5538
      ("0100110000000000", '1', '0', "--", "000", "100", "---", '1', '-', "--"), -- i=5539
      ("0100110000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5540
      ("0000010000010111", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5541
      ("0000110000010111", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5542
      ("0000110000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5543
      ("1000010000010000", '0', '1', "00", "001", "000", "100", '0', '-', "00"), -- i=5544
      ("1000110000010000", '1', '1', "00", "001", "000", "100", '0', '-', "00"), -- i=5545
      ("1000110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5546
      ("1001010000010000", '0', '1', "01", "001", "000", "100", '0', '-', "00"), -- i=5547
      ("1001110000010000", '1', '1', "01", "001", "000", "100", '0', '-', "00"), -- i=5548
      ("1001110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5549
      ("1010010000010000", '0', '1', "10", "001", "000", "100", '0', '-', "00"), -- i=5550
      ("1010110000010000", '1', '1', "10", "001", "000", "100", '0', '-', "00"), -- i=5551
      ("1010110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5552
      ("1011010000010000", '0', '1', "11", "001", "000", "100", '0', '-', "00"), -- i=5553
      ("1011110000010000", '1', '1', "11", "001", "000", "100", '0', '-', "00"), -- i=5554
      ("1011110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5555
      ("0101010000010000", '0', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5556
      ("0101110000010000", '1', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5557
      ("0101110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5558
      ("0100010000010000", '0', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5559
      ("0100110000010000", '1', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5560
      ("0100110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5561
      ("0000010011110110", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5562
      ("0000110011110110", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5563
      ("0000110011110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5564
      ("1000010000010001", '0', '1', "00", "001", "001", "100", '0', '-', "00"), -- i=5565
      ("1000110000010001", '1', '1', "00", "001", "001", "100", '0', '-', "00"), -- i=5566
      ("1000110000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5567
      ("1001010000010001", '0', '1', "01", "001", "001", "100", '0', '-', "00"), -- i=5568
      ("1001110000010001", '1', '1', "01", "001", "001", "100", '0', '-', "00"), -- i=5569
      ("1001110000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5570
      ("1010010000010001", '0', '1', "10", "001", "001", "100", '0', '-', "00"), -- i=5571
      ("1010110000010001", '1', '1', "10", "001", "001", "100", '0', '-', "00"), -- i=5572
      ("1010110000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5573
      ("1011010000010001", '0', '1', "11", "001", "001", "100", '0', '-', "00"), -- i=5574
      ("1011110000010001", '1', '1', "11", "001", "001", "100", '0', '-', "00"), -- i=5575
      ("1011110000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5576
      ("0101010000010000", '0', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5577
      ("0101110000010000", '1', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5578
      ("0101110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5579
      ("0100010000010000", '0', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5580
      ("0100110000010000", '1', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5581
      ("0100110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5582
      ("0000010010111101", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5583
      ("0000110010111101", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5584
      ("0000110010111101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5585
      ("1000010000010010", '0', '1', "00", "001", "010", "100", '0', '-', "00"), -- i=5586
      ("1000110000010010", '1', '1', "00", "001", "010", "100", '0', '-', "00"), -- i=5587
      ("1000110000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5588
      ("1001010000010010", '0', '1', "01", "001", "010", "100", '0', '-', "00"), -- i=5589
      ("1001110000010010", '1', '1', "01", "001", "010", "100", '0', '-', "00"), -- i=5590
      ("1001110000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5591
      ("1010010000010010", '0', '1', "10", "001", "010", "100", '0', '-', "00"), -- i=5592
      ("1010110000010010", '1', '1', "10", "001", "010", "100", '0', '-', "00"), -- i=5593
      ("1010110000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5594
      ("1011010000010010", '0', '1', "11", "001", "010", "100", '0', '-', "00"), -- i=5595
      ("1011110000010010", '1', '1', "11", "001", "010", "100", '0', '-', "00"), -- i=5596
      ("1011110000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5597
      ("0101010000010000", '0', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5598
      ("0101110000010000", '1', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5599
      ("0101110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5600
      ("0100010000010000", '0', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5601
      ("0100110000010000", '1', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5602
      ("0100110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5603
      ("0000010010000111", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5604
      ("0000110010000111", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5605
      ("0000110010000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5606
      ("1000010000010011", '0', '1', "00", "001", "011", "100", '0', '-', "00"), -- i=5607
      ("1000110000010011", '1', '1', "00", "001", "011", "100", '0', '-', "00"), -- i=5608
      ("1000110000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5609
      ("1001010000010011", '0', '1', "01", "001", "011", "100", '0', '-', "00"), -- i=5610
      ("1001110000010011", '1', '1', "01", "001", "011", "100", '0', '-', "00"), -- i=5611
      ("1001110000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5612
      ("1010010000010011", '0', '1', "10", "001", "011", "100", '0', '-', "00"), -- i=5613
      ("1010110000010011", '1', '1', "10", "001", "011", "100", '0', '-', "00"), -- i=5614
      ("1010110000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5615
      ("1011010000010011", '0', '1', "11", "001", "011", "100", '0', '-', "00"), -- i=5616
      ("1011110000010011", '1', '1', "11", "001", "011", "100", '0', '-', "00"), -- i=5617
      ("1011110000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5618
      ("0101010000010000", '0', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5619
      ("0101110000010000", '1', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5620
      ("0101110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5621
      ("0100010000010000", '0', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5622
      ("0100110000010000", '1', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5623
      ("0100110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5624
      ("0000010001100110", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5625
      ("0000110001100110", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5626
      ("0000110001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5627
      ("1000010000010100", '0', '1', "00", "001", "100", "100", '0', '-', "00"), -- i=5628
      ("1000110000010100", '1', '1', "00", "001", "100", "100", '0', '-', "00"), -- i=5629
      ("1000110000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5630
      ("1001010000010100", '0', '1', "01", "001", "100", "100", '0', '-', "00"), -- i=5631
      ("1001110000010100", '1', '1', "01", "001", "100", "100", '0', '-', "00"), -- i=5632
      ("1001110000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5633
      ("1010010000010100", '0', '1', "10", "001", "100", "100", '0', '-', "00"), -- i=5634
      ("1010110000010100", '1', '1', "10", "001", "100", "100", '0', '-', "00"), -- i=5635
      ("1010110000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5636
      ("1011010000010100", '0', '1', "11", "001", "100", "100", '0', '-', "00"), -- i=5637
      ("1011110000010100", '1', '1', "11", "001", "100", "100", '0', '-', "00"), -- i=5638
      ("1011110000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5639
      ("0101010000010000", '0', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5640
      ("0101110000010000", '1', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5641
      ("0101110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5642
      ("0100010000010000", '0', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5643
      ("0100110000010000", '1', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5644
      ("0100110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5645
      ("0000010000101000", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5646
      ("0000110000101000", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5647
      ("0000110000101000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5648
      ("1000010000010101", '0', '1', "00", "001", "101", "100", '0', '-', "00"), -- i=5649
      ("1000110000010101", '1', '1', "00", "001", "101", "100", '0', '-', "00"), -- i=5650
      ("1000110000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5651
      ("1001010000010101", '0', '1', "01", "001", "101", "100", '0', '-', "00"), -- i=5652
      ("1001110000010101", '1', '1', "01", "001", "101", "100", '0', '-', "00"), -- i=5653
      ("1001110000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5654
      ("1010010000010101", '0', '1', "10", "001", "101", "100", '0', '-', "00"), -- i=5655
      ("1010110000010101", '1', '1', "10", "001", "101", "100", '0', '-', "00"), -- i=5656
      ("1010110000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5657
      ("1011010000010101", '0', '1', "11", "001", "101", "100", '0', '-', "00"), -- i=5658
      ("1011110000010101", '1', '1', "11", "001", "101", "100", '0', '-', "00"), -- i=5659
      ("1011110000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5660
      ("0101010000010000", '0', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5661
      ("0101110000010000", '1', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5662
      ("0101110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5663
      ("0100010000010000", '0', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5664
      ("0100110000010000", '1', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5665
      ("0100110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5666
      ("0000010001100010", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5667
      ("0000110001100010", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5668
      ("0000110001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5669
      ("1000010000010110", '0', '1', "00", "001", "110", "100", '0', '-', "00"), -- i=5670
      ("1000110000010110", '1', '1', "00", "001", "110", "100", '0', '-', "00"), -- i=5671
      ("1000110000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5672
      ("1001010000010110", '0', '1', "01", "001", "110", "100", '0', '-', "00"), -- i=5673
      ("1001110000010110", '1', '1', "01", "001", "110", "100", '0', '-', "00"), -- i=5674
      ("1001110000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5675
      ("1010010000010110", '0', '1', "10", "001", "110", "100", '0', '-', "00"), -- i=5676
      ("1010110000010110", '1', '1', "10", "001", "110", "100", '0', '-', "00"), -- i=5677
      ("1010110000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5678
      ("1011010000010110", '0', '1', "11", "001", "110", "100", '0', '-', "00"), -- i=5679
      ("1011110000010110", '1', '1', "11", "001", "110", "100", '0', '-', "00"), -- i=5680
      ("1011110000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5681
      ("0101010000010000", '0', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5682
      ("0101110000010000", '1', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5683
      ("0101110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5684
      ("0100010000010000", '0', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5685
      ("0100110000010000", '1', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5686
      ("0100110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5687
      ("0000010011100001", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5688
      ("0000110011100001", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5689
      ("0000110011100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5690
      ("1000010000010111", '0', '1', "00", "001", "111", "100", '0', '-', "00"), -- i=5691
      ("1000110000010111", '1', '1', "00", "001", "111", "100", '0', '-', "00"), -- i=5692
      ("1000110000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5693
      ("1001010000010111", '0', '1', "01", "001", "111", "100", '0', '-', "00"), -- i=5694
      ("1001110000010111", '1', '1', "01", "001", "111", "100", '0', '-', "00"), -- i=5695
      ("1001110000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5696
      ("1010010000010111", '0', '1', "10", "001", "111", "100", '0', '-', "00"), -- i=5697
      ("1010110000010111", '1', '1', "10", "001", "111", "100", '0', '-', "00"), -- i=5698
      ("1010110000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5699
      ("1011010000010111", '0', '1', "11", "001", "111", "100", '0', '-', "00"), -- i=5700
      ("1011110000010111", '1', '1', "11", "001", "111", "100", '0', '-', "00"), -- i=5701
      ("1011110000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5702
      ("0101010000010000", '0', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5703
      ("0101110000010000", '1', '1', "--", "001", "---", "100", '0', '1', "01"), -- i=5704
      ("0101110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5705
      ("0100010000010000", '0', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5706
      ("0100110000010000", '1', '0', "--", "001", "100", "---", '1', '-', "--"), -- i=5707
      ("0100110000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5708
      ("0000010011011110", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5709
      ("0000110011011110", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5710
      ("0000110011011110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5711
      ("1000010000100000", '0', '1', "00", "010", "000", "100", '0', '-', "00"), -- i=5712
      ("1000110000100000", '1', '1', "00", "010", "000", "100", '0', '-', "00"), -- i=5713
      ("1000110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5714
      ("1001010000100000", '0', '1', "01", "010", "000", "100", '0', '-', "00"), -- i=5715
      ("1001110000100000", '1', '1', "01", "010", "000", "100", '0', '-', "00"), -- i=5716
      ("1001110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5717
      ("1010010000100000", '0', '1', "10", "010", "000", "100", '0', '-', "00"), -- i=5718
      ("1010110000100000", '1', '1', "10", "010", "000", "100", '0', '-', "00"), -- i=5719
      ("1010110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5720
      ("1011010000100000", '0', '1', "11", "010", "000", "100", '0', '-', "00"), -- i=5721
      ("1011110000100000", '1', '1', "11", "010", "000", "100", '0', '-', "00"), -- i=5722
      ("1011110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5723
      ("0101010000100000", '0', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5724
      ("0101110000100000", '1', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5725
      ("0101110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5726
      ("0100010000100000", '0', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5727
      ("0100110000100000", '1', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5728
      ("0100110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5729
      ("0000010001000110", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5730
      ("0000110001000110", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5731
      ("0000110001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5732
      ("1000010000100001", '0', '1', "00", "010", "001", "100", '0', '-', "00"), -- i=5733
      ("1000110000100001", '1', '1', "00", "010", "001", "100", '0', '-', "00"), -- i=5734
      ("1000110000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5735
      ("1001010000100001", '0', '1', "01", "010", "001", "100", '0', '-', "00"), -- i=5736
      ("1001110000100001", '1', '1', "01", "010", "001", "100", '0', '-', "00"), -- i=5737
      ("1001110000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5738
      ("1010010000100001", '0', '1', "10", "010", "001", "100", '0', '-', "00"), -- i=5739
      ("1010110000100001", '1', '1', "10", "010", "001", "100", '0', '-', "00"), -- i=5740
      ("1010110000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5741
      ("1011010000100001", '0', '1', "11", "010", "001", "100", '0', '-', "00"), -- i=5742
      ("1011110000100001", '1', '1', "11", "010", "001", "100", '0', '-', "00"), -- i=5743
      ("1011110000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5744
      ("0101010000100000", '0', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5745
      ("0101110000100000", '1', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5746
      ("0101110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5747
      ("0100010000100000", '0', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5748
      ("0100110000100000", '1', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5749
      ("0100110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5750
      ("0000010000110011", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5751
      ("0000110000110011", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5752
      ("0000110000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5753
      ("1000010000100010", '0', '1', "00", "010", "010", "100", '0', '-', "00"), -- i=5754
      ("1000110000100010", '1', '1', "00", "010", "010", "100", '0', '-', "00"), -- i=5755
      ("1000110000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5756
      ("1001010000100010", '0', '1', "01", "010", "010", "100", '0', '-', "00"), -- i=5757
      ("1001110000100010", '1', '1', "01", "010", "010", "100", '0', '-', "00"), -- i=5758
      ("1001110000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5759
      ("1010010000100010", '0', '1', "10", "010", "010", "100", '0', '-', "00"), -- i=5760
      ("1010110000100010", '1', '1', "10", "010", "010", "100", '0', '-', "00"), -- i=5761
      ("1010110000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5762
      ("1011010000100010", '0', '1', "11", "010", "010", "100", '0', '-', "00"), -- i=5763
      ("1011110000100010", '1', '1', "11", "010", "010", "100", '0', '-', "00"), -- i=5764
      ("1011110000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5765
      ("0101010000100000", '0', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5766
      ("0101110000100000", '1', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5767
      ("0101110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5768
      ("0100010000100000", '0', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5769
      ("0100110000100000", '1', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5770
      ("0100110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5771
      ("0000010000000101", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5772
      ("0000110000000101", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5773
      ("0000110000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5774
      ("1000010000100011", '0', '1', "00", "010", "011", "100", '0', '-', "00"), -- i=5775
      ("1000110000100011", '1', '1', "00", "010", "011", "100", '0', '-', "00"), -- i=5776
      ("1000110000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5777
      ("1001010000100011", '0', '1', "01", "010", "011", "100", '0', '-', "00"), -- i=5778
      ("1001110000100011", '1', '1', "01", "010", "011", "100", '0', '-', "00"), -- i=5779
      ("1001110000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5780
      ("1010010000100011", '0', '1', "10", "010", "011", "100", '0', '-', "00"), -- i=5781
      ("1010110000100011", '1', '1', "10", "010", "011", "100", '0', '-', "00"), -- i=5782
      ("1010110000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5783
      ("1011010000100011", '0', '1', "11", "010", "011", "100", '0', '-', "00"), -- i=5784
      ("1011110000100011", '1', '1', "11", "010", "011", "100", '0', '-', "00"), -- i=5785
      ("1011110000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5786
      ("0101010000100000", '0', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5787
      ("0101110000100000", '1', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5788
      ("0101110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5789
      ("0100010000100000", '0', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5790
      ("0100110000100000", '1', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5791
      ("0100110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5792
      ("0000010000111001", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5793
      ("0000110000111001", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5794
      ("0000110000111001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5795
      ("1000010000100100", '0', '1', "00", "010", "100", "100", '0', '-', "00"), -- i=5796
      ("1000110000100100", '1', '1', "00", "010", "100", "100", '0', '-', "00"), -- i=5797
      ("1000110000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5798
      ("1001010000100100", '0', '1', "01", "010", "100", "100", '0', '-', "00"), -- i=5799
      ("1001110000100100", '1', '1', "01", "010", "100", "100", '0', '-', "00"), -- i=5800
      ("1001110000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5801
      ("1010010000100100", '0', '1', "10", "010", "100", "100", '0', '-', "00"), -- i=5802
      ("1010110000100100", '1', '1', "10", "010", "100", "100", '0', '-', "00"), -- i=5803
      ("1010110000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5804
      ("1011010000100100", '0', '1', "11", "010", "100", "100", '0', '-', "00"), -- i=5805
      ("1011110000100100", '1', '1', "11", "010", "100", "100", '0', '-', "00"), -- i=5806
      ("1011110000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5807
      ("0101010000100000", '0', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5808
      ("0101110000100000", '1', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5809
      ("0101110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5810
      ("0100010000100000", '0', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5811
      ("0100110000100000", '1', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5812
      ("0100110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5813
      ("0000010001101001", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5814
      ("0000110001101001", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5815
      ("0000110001101001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5816
      ("1000010000100101", '0', '1', "00", "010", "101", "100", '0', '-', "00"), -- i=5817
      ("1000110000100101", '1', '1', "00", "010", "101", "100", '0', '-', "00"), -- i=5818
      ("1000110000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5819
      ("1001010000100101", '0', '1', "01", "010", "101", "100", '0', '-', "00"), -- i=5820
      ("1001110000100101", '1', '1', "01", "010", "101", "100", '0', '-', "00"), -- i=5821
      ("1001110000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5822
      ("1010010000100101", '0', '1', "10", "010", "101", "100", '0', '-', "00"), -- i=5823
      ("1010110000100101", '1', '1', "10", "010", "101", "100", '0', '-', "00"), -- i=5824
      ("1010110000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5825
      ("1011010000100101", '0', '1', "11", "010", "101", "100", '0', '-', "00"), -- i=5826
      ("1011110000100101", '1', '1', "11", "010", "101", "100", '0', '-', "00"), -- i=5827
      ("1011110000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5828
      ("0101010000100000", '0', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5829
      ("0101110000100000", '1', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5830
      ("0101110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5831
      ("0100010000100000", '0', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5832
      ("0100110000100000", '1', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5833
      ("0100110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5834
      ("0000010011011110", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5835
      ("0000110011011110", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5836
      ("0000110011011110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5837
      ("1000010000100110", '0', '1', "00", "010", "110", "100", '0', '-', "00"), -- i=5838
      ("1000110000100110", '1', '1', "00", "010", "110", "100", '0', '-', "00"), -- i=5839
      ("1000110000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5840
      ("1001010000100110", '0', '1', "01", "010", "110", "100", '0', '-', "00"), -- i=5841
      ("1001110000100110", '1', '1', "01", "010", "110", "100", '0', '-', "00"), -- i=5842
      ("1001110000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5843
      ("1010010000100110", '0', '1', "10", "010", "110", "100", '0', '-', "00"), -- i=5844
      ("1010110000100110", '1', '1', "10", "010", "110", "100", '0', '-', "00"), -- i=5845
      ("1010110000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5846
      ("1011010000100110", '0', '1', "11", "010", "110", "100", '0', '-', "00"), -- i=5847
      ("1011110000100110", '1', '1', "11", "010", "110", "100", '0', '-', "00"), -- i=5848
      ("1011110000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5849
      ("0101010000100000", '0', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5850
      ("0101110000100000", '1', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5851
      ("0101110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5852
      ("0100010000100000", '0', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5853
      ("0100110000100000", '1', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5854
      ("0100110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5855
      ("0000010011101001", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5856
      ("0000110011101001", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5857
      ("0000110011101001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5858
      ("1000010000100111", '0', '1', "00", "010", "111", "100", '0', '-', "00"), -- i=5859
      ("1000110000100111", '1', '1', "00", "010", "111", "100", '0', '-', "00"), -- i=5860
      ("1000110000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5861
      ("1001010000100111", '0', '1', "01", "010", "111", "100", '0', '-', "00"), -- i=5862
      ("1001110000100111", '1', '1', "01", "010", "111", "100", '0', '-', "00"), -- i=5863
      ("1001110000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5864
      ("1010010000100111", '0', '1', "10", "010", "111", "100", '0', '-', "00"), -- i=5865
      ("1010110000100111", '1', '1', "10", "010", "111", "100", '0', '-', "00"), -- i=5866
      ("1010110000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5867
      ("1011010000100111", '0', '1', "11", "010", "111", "100", '0', '-', "00"), -- i=5868
      ("1011110000100111", '1', '1', "11", "010", "111", "100", '0', '-', "00"), -- i=5869
      ("1011110000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5870
      ("0101010000100000", '0', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5871
      ("0101110000100000", '1', '1', "--", "010", "---", "100", '0', '1', "01"), -- i=5872
      ("0101110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5873
      ("0100010000100000", '0', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5874
      ("0100110000100000", '1', '0', "--", "010", "100", "---", '1', '-', "--"), -- i=5875
      ("0100110000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5876
      ("0000010011001001", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5877
      ("0000110011001001", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5878
      ("0000110011001001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5879
      ("1000010000110000", '0', '1', "00", "011", "000", "100", '0', '-', "00"), -- i=5880
      ("1000110000110000", '1', '1', "00", "011", "000", "100", '0', '-', "00"), -- i=5881
      ("1000110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5882
      ("1001010000110000", '0', '1', "01", "011", "000", "100", '0', '-', "00"), -- i=5883
      ("1001110000110000", '1', '1', "01", "011", "000", "100", '0', '-', "00"), -- i=5884
      ("1001110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5885
      ("1010010000110000", '0', '1', "10", "011", "000", "100", '0', '-', "00"), -- i=5886
      ("1010110000110000", '1', '1', "10", "011", "000", "100", '0', '-', "00"), -- i=5887
      ("1010110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5888
      ("1011010000110000", '0', '1', "11", "011", "000", "100", '0', '-', "00"), -- i=5889
      ("1011110000110000", '1', '1', "11", "011", "000", "100", '0', '-', "00"), -- i=5890
      ("1011110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5891
      ("0101010000110000", '0', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=5892
      ("0101110000110000", '1', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=5893
      ("0101110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5894
      ("0100010000110000", '0', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=5895
      ("0100110000110000", '1', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=5896
      ("0100110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5897
      ("0000010001110111", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5898
      ("0000110001110111", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5899
      ("0000110001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5900
      ("1000010000110001", '0', '1', "00", "011", "001", "100", '0', '-', "00"), -- i=5901
      ("1000110000110001", '1', '1', "00", "011", "001", "100", '0', '-', "00"), -- i=5902
      ("1000110000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5903
      ("1001010000110001", '0', '1', "01", "011", "001", "100", '0', '-', "00"), -- i=5904
      ("1001110000110001", '1', '1', "01", "011", "001", "100", '0', '-', "00"), -- i=5905
      ("1001110000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5906
      ("1010010000110001", '0', '1', "10", "011", "001", "100", '0', '-', "00"), -- i=5907
      ("1010110000110001", '1', '1', "10", "011", "001", "100", '0', '-', "00"), -- i=5908
      ("1010110000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5909
      ("1011010000110001", '0', '1', "11", "011", "001", "100", '0', '-', "00"), -- i=5910
      ("1011110000110001", '1', '1', "11", "011", "001", "100", '0', '-', "00"), -- i=5911
      ("1011110000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5912
      ("0101010000110000", '0', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=5913
      ("0101110000110000", '1', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=5914
      ("0101110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5915
      ("0100010000110000", '0', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=5916
      ("0100110000110000", '1', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=5917
      ("0100110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5918
      ("0000010011101011", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5919
      ("0000110011101011", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5920
      ("0000110011101011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5921
      ("1000010000110010", '0', '1', "00", "011", "010", "100", '0', '-', "00"), -- i=5922
      ("1000110000110010", '1', '1', "00", "011", "010", "100", '0', '-', "00"), -- i=5923
      ("1000110000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5924
      ("1001010000110010", '0', '1', "01", "011", "010", "100", '0', '-', "00"), -- i=5925
      ("1001110000110010", '1', '1', "01", "011", "010", "100", '0', '-', "00"), -- i=5926
      ("1001110000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5927
      ("1010010000110010", '0', '1', "10", "011", "010", "100", '0', '-', "00"), -- i=5928
      ("1010110000110010", '1', '1', "10", "011", "010", "100", '0', '-', "00"), -- i=5929
      ("1010110000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5930
      ("1011010000110010", '0', '1', "11", "011", "010", "100", '0', '-', "00"), -- i=5931
      ("1011110000110010", '1', '1', "11", "011", "010", "100", '0', '-', "00"), -- i=5932
      ("1011110000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5933
      ("0101010000110000", '0', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=5934
      ("0101110000110000", '1', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=5935
      ("0101110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5936
      ("0100010000110000", '0', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=5937
      ("0100110000110000", '1', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=5938
      ("0100110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5939
      ("0000010010101001", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5940
      ("0000110010101001", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5941
      ("0000110010101001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5942
      ("1000010000110011", '0', '1', "00", "011", "011", "100", '0', '-', "00"), -- i=5943
      ("1000110000110011", '1', '1', "00", "011", "011", "100", '0', '-', "00"), -- i=5944
      ("1000110000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5945
      ("1001010000110011", '0', '1', "01", "011", "011", "100", '0', '-', "00"), -- i=5946
      ("1001110000110011", '1', '1', "01", "011", "011", "100", '0', '-', "00"), -- i=5947
      ("1001110000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5948
      ("1010010000110011", '0', '1', "10", "011", "011", "100", '0', '-', "00"), -- i=5949
      ("1010110000110011", '1', '1', "10", "011", "011", "100", '0', '-', "00"), -- i=5950
      ("1010110000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5951
      ("1011010000110011", '0', '1', "11", "011", "011", "100", '0', '-', "00"), -- i=5952
      ("1011110000110011", '1', '1', "11", "011", "011", "100", '0', '-', "00"), -- i=5953
      ("1011110000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5954
      ("0101010000110000", '0', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=5955
      ("0101110000110000", '1', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=5956
      ("0101110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5957
      ("0100010000110000", '0', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=5958
      ("0100110000110000", '1', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=5959
      ("0100110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5960
      ("0000010010110111", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5961
      ("0000110010110111", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5962
      ("0000110010110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5963
      ("1000010000110100", '0', '1', "00", "011", "100", "100", '0', '-', "00"), -- i=5964
      ("1000110000110100", '1', '1', "00", "011", "100", "100", '0', '-', "00"), -- i=5965
      ("1000110000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5966
      ("1001010000110100", '0', '1', "01", "011", "100", "100", '0', '-', "00"), -- i=5967
      ("1001110000110100", '1', '1', "01", "011", "100", "100", '0', '-', "00"), -- i=5968
      ("1001110000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5969
      ("1010010000110100", '0', '1', "10", "011", "100", "100", '0', '-', "00"), -- i=5970
      ("1010110000110100", '1', '1', "10", "011", "100", "100", '0', '-', "00"), -- i=5971
      ("1010110000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5972
      ("1011010000110100", '0', '1', "11", "011", "100", "100", '0', '-', "00"), -- i=5973
      ("1011110000110100", '1', '1', "11", "011", "100", "100", '0', '-', "00"), -- i=5974
      ("1011110000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5975
      ("0101010000110000", '0', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=5976
      ("0101110000110000", '1', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=5977
      ("0101110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5978
      ("0100010000110000", '0', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=5979
      ("0100110000110000", '1', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=5980
      ("0100110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5981
      ("0000010011111000", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5982
      ("0000110011111000", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=5983
      ("0000110011111000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5984
      ("1000010000110101", '0', '1', "00", "011", "101", "100", '0', '-', "00"), -- i=5985
      ("1000110000110101", '1', '1', "00", "011", "101", "100", '0', '-', "00"), -- i=5986
      ("1000110000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5987
      ("1001010000110101", '0', '1', "01", "011", "101", "100", '0', '-', "00"), -- i=5988
      ("1001110000110101", '1', '1', "01", "011", "101", "100", '0', '-', "00"), -- i=5989
      ("1001110000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5990
      ("1010010000110101", '0', '1', "10", "011", "101", "100", '0', '-', "00"), -- i=5991
      ("1010110000110101", '1', '1', "10", "011", "101", "100", '0', '-', "00"), -- i=5992
      ("1010110000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5993
      ("1011010000110101", '0', '1', "11", "011", "101", "100", '0', '-', "00"), -- i=5994
      ("1011110000110101", '1', '1', "11", "011", "101", "100", '0', '-', "00"), -- i=5995
      ("1011110000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5996
      ("0101010000110000", '0', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=5997
      ("0101110000110000", '1', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=5998
      ("0101110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=5999
      ("0100010000110000", '0', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=6000
      ("0100110000110000", '1', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=6001
      ("0100110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6002
      ("0000010010111011", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6003
      ("0000110010111011", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6004
      ("0000110010111011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6005
      ("1000010000110110", '0', '1', "00", "011", "110", "100", '0', '-', "00"), -- i=6006
      ("1000110000110110", '1', '1', "00", "011", "110", "100", '0', '-', "00"), -- i=6007
      ("1000110000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6008
      ("1001010000110110", '0', '1', "01", "011", "110", "100", '0', '-', "00"), -- i=6009
      ("1001110000110110", '1', '1', "01", "011", "110", "100", '0', '-', "00"), -- i=6010
      ("1001110000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6011
      ("1010010000110110", '0', '1', "10", "011", "110", "100", '0', '-', "00"), -- i=6012
      ("1010110000110110", '1', '1', "10", "011", "110", "100", '0', '-', "00"), -- i=6013
      ("1010110000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6014
      ("1011010000110110", '0', '1', "11", "011", "110", "100", '0', '-', "00"), -- i=6015
      ("1011110000110110", '1', '1', "11", "011", "110", "100", '0', '-', "00"), -- i=6016
      ("1011110000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6017
      ("0101010000110000", '0', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=6018
      ("0101110000110000", '1', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=6019
      ("0101110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6020
      ("0100010000110000", '0', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=6021
      ("0100110000110000", '1', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=6022
      ("0100110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6023
      ("0000010000100101", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6024
      ("0000110000100101", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6025
      ("0000110000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6026
      ("1000010000110111", '0', '1', "00", "011", "111", "100", '0', '-', "00"), -- i=6027
      ("1000110000110111", '1', '1', "00", "011", "111", "100", '0', '-', "00"), -- i=6028
      ("1000110000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6029
      ("1001010000110111", '0', '1', "01", "011", "111", "100", '0', '-', "00"), -- i=6030
      ("1001110000110111", '1', '1', "01", "011", "111", "100", '0', '-', "00"), -- i=6031
      ("1001110000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6032
      ("1010010000110111", '0', '1', "10", "011", "111", "100", '0', '-', "00"), -- i=6033
      ("1010110000110111", '1', '1', "10", "011", "111", "100", '0', '-', "00"), -- i=6034
      ("1010110000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6035
      ("1011010000110111", '0', '1', "11", "011", "111", "100", '0', '-', "00"), -- i=6036
      ("1011110000110111", '1', '1', "11", "011", "111", "100", '0', '-', "00"), -- i=6037
      ("1011110000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6038
      ("0101010000110000", '0', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=6039
      ("0101110000110000", '1', '1', "--", "011", "---", "100", '0', '1', "01"), -- i=6040
      ("0101110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6041
      ("0100010000110000", '0', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=6042
      ("0100110000110000", '1', '0', "--", "011", "100", "---", '1', '-', "--"), -- i=6043
      ("0100110000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6044
      ("0000010001001100", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6045
      ("0000110001001100", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6046
      ("0000110001001100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6047
      ("1000010001000000", '0', '1', "00", "100", "000", "100", '0', '-', "00"), -- i=6048
      ("1000110001000000", '1', '1', "00", "100", "000", "100", '0', '-', "00"), -- i=6049
      ("1000110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6050
      ("1001010001000000", '0', '1', "01", "100", "000", "100", '0', '-', "00"), -- i=6051
      ("1001110001000000", '1', '1', "01", "100", "000", "100", '0', '-', "00"), -- i=6052
      ("1001110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6053
      ("1010010001000000", '0', '1', "10", "100", "000", "100", '0', '-', "00"), -- i=6054
      ("1010110001000000", '1', '1', "10", "100", "000", "100", '0', '-', "00"), -- i=6055
      ("1010110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6056
      ("1011010001000000", '0', '1', "11", "100", "000", "100", '0', '-', "00"), -- i=6057
      ("1011110001000000", '1', '1', "11", "100", "000", "100", '0', '-', "00"), -- i=6058
      ("1011110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6059
      ("0101010001000000", '0', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6060
      ("0101110001000000", '1', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6061
      ("0101110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6062
      ("0100010001000000", '0', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6063
      ("0100110001000000", '1', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6064
      ("0100110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6065
      ("0000010010101000", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6066
      ("0000110010101000", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6067
      ("0000110010101000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6068
      ("1000010001000001", '0', '1', "00", "100", "001", "100", '0', '-', "00"), -- i=6069
      ("1000110001000001", '1', '1', "00", "100", "001", "100", '0', '-', "00"), -- i=6070
      ("1000110001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6071
      ("1001010001000001", '0', '1', "01", "100", "001", "100", '0', '-', "00"), -- i=6072
      ("1001110001000001", '1', '1', "01", "100", "001", "100", '0', '-', "00"), -- i=6073
      ("1001110001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6074
      ("1010010001000001", '0', '1', "10", "100", "001", "100", '0', '-', "00"), -- i=6075
      ("1010110001000001", '1', '1', "10", "100", "001", "100", '0', '-', "00"), -- i=6076
      ("1010110001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6077
      ("1011010001000001", '0', '1', "11", "100", "001", "100", '0', '-', "00"), -- i=6078
      ("1011110001000001", '1', '1', "11", "100", "001", "100", '0', '-', "00"), -- i=6079
      ("1011110001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6080
      ("0101010001000000", '0', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6081
      ("0101110001000000", '1', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6082
      ("0101110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6083
      ("0100010001000000", '0', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6084
      ("0100110001000000", '1', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6085
      ("0100110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6086
      ("0000010001000100", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6087
      ("0000110001000100", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6088
      ("0000110001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6089
      ("1000010001000010", '0', '1', "00", "100", "010", "100", '0', '-', "00"), -- i=6090
      ("1000110001000010", '1', '1', "00", "100", "010", "100", '0', '-', "00"), -- i=6091
      ("1000110001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6092
      ("1001010001000010", '0', '1', "01", "100", "010", "100", '0', '-', "00"), -- i=6093
      ("1001110001000010", '1', '1', "01", "100", "010", "100", '0', '-', "00"), -- i=6094
      ("1001110001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6095
      ("1010010001000010", '0', '1', "10", "100", "010", "100", '0', '-', "00"), -- i=6096
      ("1010110001000010", '1', '1', "10", "100", "010", "100", '0', '-', "00"), -- i=6097
      ("1010110001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6098
      ("1011010001000010", '0', '1', "11", "100", "010", "100", '0', '-', "00"), -- i=6099
      ("1011110001000010", '1', '1', "11", "100", "010", "100", '0', '-', "00"), -- i=6100
      ("1011110001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6101
      ("0101010001000000", '0', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6102
      ("0101110001000000", '1', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6103
      ("0101110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6104
      ("0100010001000000", '0', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6105
      ("0100110001000000", '1', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6106
      ("0100110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6107
      ("0000010000111001", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6108
      ("0000110000111001", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6109
      ("0000110000111001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6110
      ("1000010001000011", '0', '1', "00", "100", "011", "100", '0', '-', "00"), -- i=6111
      ("1000110001000011", '1', '1', "00", "100", "011", "100", '0', '-', "00"), -- i=6112
      ("1000110001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6113
      ("1001010001000011", '0', '1', "01", "100", "011", "100", '0', '-', "00"), -- i=6114
      ("1001110001000011", '1', '1', "01", "100", "011", "100", '0', '-', "00"), -- i=6115
      ("1001110001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6116
      ("1010010001000011", '0', '1', "10", "100", "011", "100", '0', '-', "00"), -- i=6117
      ("1010110001000011", '1', '1', "10", "100", "011", "100", '0', '-', "00"), -- i=6118
      ("1010110001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6119
      ("1011010001000011", '0', '1', "11", "100", "011", "100", '0', '-', "00"), -- i=6120
      ("1011110001000011", '1', '1', "11", "100", "011", "100", '0', '-', "00"), -- i=6121
      ("1011110001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6122
      ("0101010001000000", '0', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6123
      ("0101110001000000", '1', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6124
      ("0101110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6125
      ("0100010001000000", '0', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6126
      ("0100110001000000", '1', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6127
      ("0100110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6128
      ("0000010000010010", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6129
      ("0000110000010010", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6130
      ("0000110000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6131
      ("1000010001000100", '0', '1', "00", "100", "100", "100", '0', '-', "00"), -- i=6132
      ("1000110001000100", '1', '1', "00", "100", "100", "100", '0', '-', "00"), -- i=6133
      ("1000110001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6134
      ("1001010001000100", '0', '1', "01", "100", "100", "100", '0', '-', "00"), -- i=6135
      ("1001110001000100", '1', '1', "01", "100", "100", "100", '0', '-', "00"), -- i=6136
      ("1001110001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6137
      ("1010010001000100", '0', '1', "10", "100", "100", "100", '0', '-', "00"), -- i=6138
      ("1010110001000100", '1', '1', "10", "100", "100", "100", '0', '-', "00"), -- i=6139
      ("1010110001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6140
      ("1011010001000100", '0', '1', "11", "100", "100", "100", '0', '-', "00"), -- i=6141
      ("1011110001000100", '1', '1', "11", "100", "100", "100", '0', '-', "00"), -- i=6142
      ("1011110001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6143
      ("0101010001000000", '0', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6144
      ("0101110001000000", '1', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6145
      ("0101110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6146
      ("0100010001000000", '0', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6147
      ("0100110001000000", '1', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6148
      ("0100110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6149
      ("0000010000011000", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6150
      ("0000110000011000", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6151
      ("0000110000011000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6152
      ("1000010001000101", '0', '1', "00", "100", "101", "100", '0', '-', "00"), -- i=6153
      ("1000110001000101", '1', '1', "00", "100", "101", "100", '0', '-', "00"), -- i=6154
      ("1000110001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6155
      ("1001010001000101", '0', '1', "01", "100", "101", "100", '0', '-', "00"), -- i=6156
      ("1001110001000101", '1', '1', "01", "100", "101", "100", '0', '-', "00"), -- i=6157
      ("1001110001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6158
      ("1010010001000101", '0', '1', "10", "100", "101", "100", '0', '-', "00"), -- i=6159
      ("1010110001000101", '1', '1', "10", "100", "101", "100", '0', '-', "00"), -- i=6160
      ("1010110001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6161
      ("1011010001000101", '0', '1', "11", "100", "101", "100", '0', '-', "00"), -- i=6162
      ("1011110001000101", '1', '1', "11", "100", "101", "100", '0', '-', "00"), -- i=6163
      ("1011110001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6164
      ("0101010001000000", '0', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6165
      ("0101110001000000", '1', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6166
      ("0101110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6167
      ("0100010001000000", '0', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6168
      ("0100110001000000", '1', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6169
      ("0100110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6170
      ("0000010000111001", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6171
      ("0000110000111001", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6172
      ("0000110000111001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6173
      ("1000010001000110", '0', '1', "00", "100", "110", "100", '0', '-', "00"), -- i=6174
      ("1000110001000110", '1', '1', "00", "100", "110", "100", '0', '-', "00"), -- i=6175
      ("1000110001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6176
      ("1001010001000110", '0', '1', "01", "100", "110", "100", '0', '-', "00"), -- i=6177
      ("1001110001000110", '1', '1', "01", "100", "110", "100", '0', '-', "00"), -- i=6178
      ("1001110001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6179
      ("1010010001000110", '0', '1', "10", "100", "110", "100", '0', '-', "00"), -- i=6180
      ("1010110001000110", '1', '1', "10", "100", "110", "100", '0', '-', "00"), -- i=6181
      ("1010110001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6182
      ("1011010001000110", '0', '1', "11", "100", "110", "100", '0', '-', "00"), -- i=6183
      ("1011110001000110", '1', '1', "11", "100", "110", "100", '0', '-', "00"), -- i=6184
      ("1011110001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6185
      ("0101010001000000", '0', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6186
      ("0101110001000000", '1', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6187
      ("0101110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6188
      ("0100010001000000", '0', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6189
      ("0100110001000000", '1', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6190
      ("0100110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6191
      ("0000010010101010", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6192
      ("0000110010101010", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6193
      ("0000110010101010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6194
      ("1000010001000111", '0', '1', "00", "100", "111", "100", '0', '-', "00"), -- i=6195
      ("1000110001000111", '1', '1', "00", "100", "111", "100", '0', '-', "00"), -- i=6196
      ("1000110001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6197
      ("1001010001000111", '0', '1', "01", "100", "111", "100", '0', '-', "00"), -- i=6198
      ("1001110001000111", '1', '1', "01", "100", "111", "100", '0', '-', "00"), -- i=6199
      ("1001110001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6200
      ("1010010001000111", '0', '1', "10", "100", "111", "100", '0', '-', "00"), -- i=6201
      ("1010110001000111", '1', '1', "10", "100", "111", "100", '0', '-', "00"), -- i=6202
      ("1010110001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6203
      ("1011010001000111", '0', '1', "11", "100", "111", "100", '0', '-', "00"), -- i=6204
      ("1011110001000111", '1', '1', "11", "100", "111", "100", '0', '-', "00"), -- i=6205
      ("1011110001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6206
      ("0101010001000000", '0', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6207
      ("0101110001000000", '1', '1', "--", "100", "---", "100", '0', '1', "01"), -- i=6208
      ("0101110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6209
      ("0100010001000000", '0', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6210
      ("0100110001000000", '1', '0', "--", "100", "100", "---", '1', '-', "--"), -- i=6211
      ("0100110001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6212
      ("0000010000100101", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6213
      ("0000110000100101", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6214
      ("0000110000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6215
      ("1000010001010000", '0', '1', "00", "101", "000", "100", '0', '-', "00"), -- i=6216
      ("1000110001010000", '1', '1', "00", "101", "000", "100", '0', '-', "00"), -- i=6217
      ("1000110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6218
      ("1001010001010000", '0', '1', "01", "101", "000", "100", '0', '-', "00"), -- i=6219
      ("1001110001010000", '1', '1', "01", "101", "000", "100", '0', '-', "00"), -- i=6220
      ("1001110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6221
      ("1010010001010000", '0', '1', "10", "101", "000", "100", '0', '-', "00"), -- i=6222
      ("1010110001010000", '1', '1', "10", "101", "000", "100", '0', '-', "00"), -- i=6223
      ("1010110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6224
      ("1011010001010000", '0', '1', "11", "101", "000", "100", '0', '-', "00"), -- i=6225
      ("1011110001010000", '1', '1', "11", "101", "000", "100", '0', '-', "00"), -- i=6226
      ("1011110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6227
      ("0101010001010000", '0', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6228
      ("0101110001010000", '1', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6229
      ("0101110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6230
      ("0100010001010000", '0', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6231
      ("0100110001010000", '1', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6232
      ("0100110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6233
      ("0000010001110100", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6234
      ("0000110001110100", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6235
      ("0000110001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6236
      ("1000010001010001", '0', '1', "00", "101", "001", "100", '0', '-', "00"), -- i=6237
      ("1000110001010001", '1', '1', "00", "101", "001", "100", '0', '-', "00"), -- i=6238
      ("1000110001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6239
      ("1001010001010001", '0', '1', "01", "101", "001", "100", '0', '-', "00"), -- i=6240
      ("1001110001010001", '1', '1', "01", "101", "001", "100", '0', '-', "00"), -- i=6241
      ("1001110001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6242
      ("1010010001010001", '0', '1', "10", "101", "001", "100", '0', '-', "00"), -- i=6243
      ("1010110001010001", '1', '1', "10", "101", "001", "100", '0', '-', "00"), -- i=6244
      ("1010110001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6245
      ("1011010001010001", '0', '1', "11", "101", "001", "100", '0', '-', "00"), -- i=6246
      ("1011110001010001", '1', '1', "11", "101", "001", "100", '0', '-', "00"), -- i=6247
      ("1011110001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6248
      ("0101010001010000", '0', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6249
      ("0101110001010000", '1', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6250
      ("0101110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6251
      ("0100010001010000", '0', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6252
      ("0100110001010000", '1', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6253
      ("0100110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6254
      ("0000010001100111", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6255
      ("0000110001100111", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6256
      ("0000110001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6257
      ("1000010001010010", '0', '1', "00", "101", "010", "100", '0', '-', "00"), -- i=6258
      ("1000110001010010", '1', '1', "00", "101", "010", "100", '0', '-', "00"), -- i=6259
      ("1000110001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6260
      ("1001010001010010", '0', '1', "01", "101", "010", "100", '0', '-', "00"), -- i=6261
      ("1001110001010010", '1', '1', "01", "101", "010", "100", '0', '-', "00"), -- i=6262
      ("1001110001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6263
      ("1010010001010010", '0', '1', "10", "101", "010", "100", '0', '-', "00"), -- i=6264
      ("1010110001010010", '1', '1', "10", "101", "010", "100", '0', '-', "00"), -- i=6265
      ("1010110001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6266
      ("1011010001010010", '0', '1', "11", "101", "010", "100", '0', '-', "00"), -- i=6267
      ("1011110001010010", '1', '1', "11", "101", "010", "100", '0', '-', "00"), -- i=6268
      ("1011110001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6269
      ("0101010001010000", '0', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6270
      ("0101110001010000", '1', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6271
      ("0101110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6272
      ("0100010001010000", '0', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6273
      ("0100110001010000", '1', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6274
      ("0100110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6275
      ("0000010001110110", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6276
      ("0000110001110110", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6277
      ("0000110001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6278
      ("1000010001010011", '0', '1', "00", "101", "011", "100", '0', '-', "00"), -- i=6279
      ("1000110001010011", '1', '1', "00", "101", "011", "100", '0', '-', "00"), -- i=6280
      ("1000110001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6281
      ("1001010001010011", '0', '1', "01", "101", "011", "100", '0', '-', "00"), -- i=6282
      ("1001110001010011", '1', '1', "01", "101", "011", "100", '0', '-', "00"), -- i=6283
      ("1001110001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6284
      ("1010010001010011", '0', '1', "10", "101", "011", "100", '0', '-', "00"), -- i=6285
      ("1010110001010011", '1', '1', "10", "101", "011", "100", '0', '-', "00"), -- i=6286
      ("1010110001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6287
      ("1011010001010011", '0', '1', "11", "101", "011", "100", '0', '-', "00"), -- i=6288
      ("1011110001010011", '1', '1', "11", "101", "011", "100", '0', '-', "00"), -- i=6289
      ("1011110001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6290
      ("0101010001010000", '0', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6291
      ("0101110001010000", '1', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6292
      ("0101110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6293
      ("0100010001010000", '0', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6294
      ("0100110001010000", '1', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6295
      ("0100110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6296
      ("0000010010110110", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6297
      ("0000110010110110", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6298
      ("0000110010110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6299
      ("1000010001010100", '0', '1', "00", "101", "100", "100", '0', '-', "00"), -- i=6300
      ("1000110001010100", '1', '1', "00", "101", "100", "100", '0', '-', "00"), -- i=6301
      ("1000110001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6302
      ("1001010001010100", '0', '1', "01", "101", "100", "100", '0', '-', "00"), -- i=6303
      ("1001110001010100", '1', '1', "01", "101", "100", "100", '0', '-', "00"), -- i=6304
      ("1001110001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6305
      ("1010010001010100", '0', '1', "10", "101", "100", "100", '0', '-', "00"), -- i=6306
      ("1010110001010100", '1', '1', "10", "101", "100", "100", '0', '-', "00"), -- i=6307
      ("1010110001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6308
      ("1011010001010100", '0', '1', "11", "101", "100", "100", '0', '-', "00"), -- i=6309
      ("1011110001010100", '1', '1', "11", "101", "100", "100", '0', '-', "00"), -- i=6310
      ("1011110001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6311
      ("0101010001010000", '0', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6312
      ("0101110001010000", '1', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6313
      ("0101110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6314
      ("0100010001010000", '0', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6315
      ("0100110001010000", '1', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6316
      ("0100110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6317
      ("0000010010101100", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6318
      ("0000110010101100", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6319
      ("0000110010101100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6320
      ("1000010001010101", '0', '1', "00", "101", "101", "100", '0', '-', "00"), -- i=6321
      ("1000110001010101", '1', '1', "00", "101", "101", "100", '0', '-', "00"), -- i=6322
      ("1000110001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6323
      ("1001010001010101", '0', '1', "01", "101", "101", "100", '0', '-', "00"), -- i=6324
      ("1001110001010101", '1', '1', "01", "101", "101", "100", '0', '-', "00"), -- i=6325
      ("1001110001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6326
      ("1010010001010101", '0', '1', "10", "101", "101", "100", '0', '-', "00"), -- i=6327
      ("1010110001010101", '1', '1', "10", "101", "101", "100", '0', '-', "00"), -- i=6328
      ("1010110001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6329
      ("1011010001010101", '0', '1', "11", "101", "101", "100", '0', '-', "00"), -- i=6330
      ("1011110001010101", '1', '1', "11", "101", "101", "100", '0', '-', "00"), -- i=6331
      ("1011110001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6332
      ("0101010001010000", '0', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6333
      ("0101110001010000", '1', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6334
      ("0101110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6335
      ("0100010001010000", '0', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6336
      ("0100110001010000", '1', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6337
      ("0100110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6338
      ("0000010010001101", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6339
      ("0000110010001101", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6340
      ("0000110010001101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6341
      ("1000010001010110", '0', '1', "00", "101", "110", "100", '0', '-', "00"), -- i=6342
      ("1000110001010110", '1', '1', "00", "101", "110", "100", '0', '-', "00"), -- i=6343
      ("1000110001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6344
      ("1001010001010110", '0', '1', "01", "101", "110", "100", '0', '-', "00"), -- i=6345
      ("1001110001010110", '1', '1', "01", "101", "110", "100", '0', '-', "00"), -- i=6346
      ("1001110001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6347
      ("1010010001010110", '0', '1', "10", "101", "110", "100", '0', '-', "00"), -- i=6348
      ("1010110001010110", '1', '1', "10", "101", "110", "100", '0', '-', "00"), -- i=6349
      ("1010110001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6350
      ("1011010001010110", '0', '1', "11", "101", "110", "100", '0', '-', "00"), -- i=6351
      ("1011110001010110", '1', '1', "11", "101", "110", "100", '0', '-', "00"), -- i=6352
      ("1011110001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6353
      ("0101010001010000", '0', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6354
      ("0101110001010000", '1', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6355
      ("0101110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6356
      ("0100010001010000", '0', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6357
      ("0100110001010000", '1', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6358
      ("0100110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6359
      ("0000010011111110", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6360
      ("0000110011111110", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6361
      ("0000110011111110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6362
      ("1000010001010111", '0', '1', "00", "101", "111", "100", '0', '-', "00"), -- i=6363
      ("1000110001010111", '1', '1', "00", "101", "111", "100", '0', '-', "00"), -- i=6364
      ("1000110001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6365
      ("1001010001010111", '0', '1', "01", "101", "111", "100", '0', '-', "00"), -- i=6366
      ("1001110001010111", '1', '1', "01", "101", "111", "100", '0', '-', "00"), -- i=6367
      ("1001110001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6368
      ("1010010001010111", '0', '1', "10", "101", "111", "100", '0', '-', "00"), -- i=6369
      ("1010110001010111", '1', '1', "10", "101", "111", "100", '0', '-', "00"), -- i=6370
      ("1010110001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6371
      ("1011010001010111", '0', '1', "11", "101", "111", "100", '0', '-', "00"), -- i=6372
      ("1011110001010111", '1', '1', "11", "101", "111", "100", '0', '-', "00"), -- i=6373
      ("1011110001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6374
      ("0101010001010000", '0', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6375
      ("0101110001010000", '1', '1', "--", "101", "---", "100", '0', '1', "01"), -- i=6376
      ("0101110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6377
      ("0100010001010000", '0', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6378
      ("0100110001010000", '1', '0', "--", "101", "100", "---", '1', '-', "--"), -- i=6379
      ("0100110001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6380
      ("0000010001011110", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6381
      ("0000110001011110", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6382
      ("0000110001011110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6383
      ("1000010001100000", '0', '1', "00", "110", "000", "100", '0', '-', "00"), -- i=6384
      ("1000110001100000", '1', '1', "00", "110", "000", "100", '0', '-', "00"), -- i=6385
      ("1000110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6386
      ("1001010001100000", '0', '1', "01", "110", "000", "100", '0', '-', "00"), -- i=6387
      ("1001110001100000", '1', '1', "01", "110", "000", "100", '0', '-', "00"), -- i=6388
      ("1001110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6389
      ("1010010001100000", '0', '1', "10", "110", "000", "100", '0', '-', "00"), -- i=6390
      ("1010110001100000", '1', '1', "10", "110", "000", "100", '0', '-', "00"), -- i=6391
      ("1010110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6392
      ("1011010001100000", '0', '1', "11", "110", "000", "100", '0', '-', "00"), -- i=6393
      ("1011110001100000", '1', '1', "11", "110", "000", "100", '0', '-', "00"), -- i=6394
      ("1011110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6395
      ("0101010001100000", '0', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6396
      ("0101110001100000", '1', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6397
      ("0101110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6398
      ("0100010001100000", '0', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6399
      ("0100110001100000", '1', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6400
      ("0100110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6401
      ("0000010001100110", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6402
      ("0000110001100110", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6403
      ("0000110001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6404
      ("1000010001100001", '0', '1', "00", "110", "001", "100", '0', '-', "00"), -- i=6405
      ("1000110001100001", '1', '1', "00", "110", "001", "100", '0', '-', "00"), -- i=6406
      ("1000110001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6407
      ("1001010001100001", '0', '1', "01", "110", "001", "100", '0', '-', "00"), -- i=6408
      ("1001110001100001", '1', '1', "01", "110", "001", "100", '0', '-', "00"), -- i=6409
      ("1001110001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6410
      ("1010010001100001", '0', '1', "10", "110", "001", "100", '0', '-', "00"), -- i=6411
      ("1010110001100001", '1', '1', "10", "110", "001", "100", '0', '-', "00"), -- i=6412
      ("1010110001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6413
      ("1011010001100001", '0', '1', "11", "110", "001", "100", '0', '-', "00"), -- i=6414
      ("1011110001100001", '1', '1', "11", "110", "001", "100", '0', '-', "00"), -- i=6415
      ("1011110001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6416
      ("0101010001100000", '0', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6417
      ("0101110001100000", '1', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6418
      ("0101110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6419
      ("0100010001100000", '0', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6420
      ("0100110001100000", '1', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6421
      ("0100110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6422
      ("0000010011100110", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6423
      ("0000110011100110", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6424
      ("0000110011100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6425
      ("1000010001100010", '0', '1', "00", "110", "010", "100", '0', '-', "00"), -- i=6426
      ("1000110001100010", '1', '1', "00", "110", "010", "100", '0', '-', "00"), -- i=6427
      ("1000110001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6428
      ("1001010001100010", '0', '1', "01", "110", "010", "100", '0', '-', "00"), -- i=6429
      ("1001110001100010", '1', '1', "01", "110", "010", "100", '0', '-', "00"), -- i=6430
      ("1001110001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6431
      ("1010010001100010", '0', '1', "10", "110", "010", "100", '0', '-', "00"), -- i=6432
      ("1010110001100010", '1', '1', "10", "110", "010", "100", '0', '-', "00"), -- i=6433
      ("1010110001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6434
      ("1011010001100010", '0', '1', "11", "110", "010", "100", '0', '-', "00"), -- i=6435
      ("1011110001100010", '1', '1', "11", "110", "010", "100", '0', '-', "00"), -- i=6436
      ("1011110001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6437
      ("0101010001100000", '0', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6438
      ("0101110001100000", '1', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6439
      ("0101110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6440
      ("0100010001100000", '0', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6441
      ("0100110001100000", '1', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6442
      ("0100110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6443
      ("0000010010101001", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6444
      ("0000110010101001", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6445
      ("0000110010101001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6446
      ("1000010001100011", '0', '1', "00", "110", "011", "100", '0', '-', "00"), -- i=6447
      ("1000110001100011", '1', '1', "00", "110", "011", "100", '0', '-', "00"), -- i=6448
      ("1000110001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6449
      ("1001010001100011", '0', '1', "01", "110", "011", "100", '0', '-', "00"), -- i=6450
      ("1001110001100011", '1', '1', "01", "110", "011", "100", '0', '-', "00"), -- i=6451
      ("1001110001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6452
      ("1010010001100011", '0', '1', "10", "110", "011", "100", '0', '-', "00"), -- i=6453
      ("1010110001100011", '1', '1', "10", "110", "011", "100", '0', '-', "00"), -- i=6454
      ("1010110001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6455
      ("1011010001100011", '0', '1', "11", "110", "011", "100", '0', '-', "00"), -- i=6456
      ("1011110001100011", '1', '1', "11", "110", "011", "100", '0', '-', "00"), -- i=6457
      ("1011110001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6458
      ("0101010001100000", '0', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6459
      ("0101110001100000", '1', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6460
      ("0101110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6461
      ("0100010001100000", '0', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6462
      ("0100110001100000", '1', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6463
      ("0100110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6464
      ("0000010010101011", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6465
      ("0000110010101011", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6466
      ("0000110010101011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6467
      ("1000010001100100", '0', '1', "00", "110", "100", "100", '0', '-', "00"), -- i=6468
      ("1000110001100100", '1', '1', "00", "110", "100", "100", '0', '-', "00"), -- i=6469
      ("1000110001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6470
      ("1001010001100100", '0', '1', "01", "110", "100", "100", '0', '-', "00"), -- i=6471
      ("1001110001100100", '1', '1', "01", "110", "100", "100", '0', '-', "00"), -- i=6472
      ("1001110001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6473
      ("1010010001100100", '0', '1', "10", "110", "100", "100", '0', '-', "00"), -- i=6474
      ("1010110001100100", '1', '1', "10", "110", "100", "100", '0', '-', "00"), -- i=6475
      ("1010110001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6476
      ("1011010001100100", '0', '1', "11", "110", "100", "100", '0', '-', "00"), -- i=6477
      ("1011110001100100", '1', '1', "11", "110", "100", "100", '0', '-', "00"), -- i=6478
      ("1011110001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6479
      ("0101010001100000", '0', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6480
      ("0101110001100000", '1', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6481
      ("0101110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6482
      ("0100010001100000", '0', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6483
      ("0100110001100000", '1', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6484
      ("0100110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6485
      ("0000010011101111", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6486
      ("0000110011101111", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6487
      ("0000110011101111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6488
      ("1000010001100101", '0', '1', "00", "110", "101", "100", '0', '-', "00"), -- i=6489
      ("1000110001100101", '1', '1', "00", "110", "101", "100", '0', '-', "00"), -- i=6490
      ("1000110001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6491
      ("1001010001100101", '0', '1', "01", "110", "101", "100", '0', '-', "00"), -- i=6492
      ("1001110001100101", '1', '1', "01", "110", "101", "100", '0', '-', "00"), -- i=6493
      ("1001110001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6494
      ("1010010001100101", '0', '1', "10", "110", "101", "100", '0', '-', "00"), -- i=6495
      ("1010110001100101", '1', '1', "10", "110", "101", "100", '0', '-', "00"), -- i=6496
      ("1010110001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6497
      ("1011010001100101", '0', '1', "11", "110", "101", "100", '0', '-', "00"), -- i=6498
      ("1011110001100101", '1', '1', "11", "110", "101", "100", '0', '-', "00"), -- i=6499
      ("1011110001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6500
      ("0101010001100000", '0', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6501
      ("0101110001100000", '1', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6502
      ("0101110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6503
      ("0100010001100000", '0', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6504
      ("0100110001100000", '1', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6505
      ("0100110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6506
      ("0000010001110100", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6507
      ("0000110001110100", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6508
      ("0000110001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6509
      ("1000010001100110", '0', '1', "00", "110", "110", "100", '0', '-', "00"), -- i=6510
      ("1000110001100110", '1', '1', "00", "110", "110", "100", '0', '-', "00"), -- i=6511
      ("1000110001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6512
      ("1001010001100110", '0', '1', "01", "110", "110", "100", '0', '-', "00"), -- i=6513
      ("1001110001100110", '1', '1', "01", "110", "110", "100", '0', '-', "00"), -- i=6514
      ("1001110001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6515
      ("1010010001100110", '0', '1', "10", "110", "110", "100", '0', '-', "00"), -- i=6516
      ("1010110001100110", '1', '1', "10", "110", "110", "100", '0', '-', "00"), -- i=6517
      ("1010110001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6518
      ("1011010001100110", '0', '1', "11", "110", "110", "100", '0', '-', "00"), -- i=6519
      ("1011110001100110", '1', '1', "11", "110", "110", "100", '0', '-', "00"), -- i=6520
      ("1011110001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6521
      ("0101010001100000", '0', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6522
      ("0101110001100000", '1', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6523
      ("0101110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6524
      ("0100010001100000", '0', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6525
      ("0100110001100000", '1', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6526
      ("0100110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6527
      ("0000010011100001", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6528
      ("0000110011100001", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6529
      ("0000110011100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6530
      ("1000010001100111", '0', '1', "00", "110", "111", "100", '0', '-', "00"), -- i=6531
      ("1000110001100111", '1', '1', "00", "110", "111", "100", '0', '-', "00"), -- i=6532
      ("1000110001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6533
      ("1001010001100111", '0', '1', "01", "110", "111", "100", '0', '-', "00"), -- i=6534
      ("1001110001100111", '1', '1', "01", "110", "111", "100", '0', '-', "00"), -- i=6535
      ("1001110001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6536
      ("1010010001100111", '0', '1', "10", "110", "111", "100", '0', '-', "00"), -- i=6537
      ("1010110001100111", '1', '1', "10", "110", "111", "100", '0', '-', "00"), -- i=6538
      ("1010110001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6539
      ("1011010001100111", '0', '1', "11", "110", "111", "100", '0', '-', "00"), -- i=6540
      ("1011110001100111", '1', '1', "11", "110", "111", "100", '0', '-', "00"), -- i=6541
      ("1011110001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6542
      ("0101010001100000", '0', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6543
      ("0101110001100000", '1', '1', "--", "110", "---", "100", '0', '1', "01"), -- i=6544
      ("0101110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6545
      ("0100010001100000", '0', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6546
      ("0100110001100000", '1', '0', "--", "110", "100", "---", '1', '-', "--"), -- i=6547
      ("0100110001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6548
      ("0000010011110011", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6549
      ("0000110011110011", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6550
      ("0000110011110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6551
      ("1000010001110000", '0', '1', "00", "111", "000", "100", '0', '-', "00"), -- i=6552
      ("1000110001110000", '1', '1', "00", "111", "000", "100", '0', '-', "00"), -- i=6553
      ("1000110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6554
      ("1001010001110000", '0', '1', "01", "111", "000", "100", '0', '-', "00"), -- i=6555
      ("1001110001110000", '1', '1', "01", "111", "000", "100", '0', '-', "00"), -- i=6556
      ("1001110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6557
      ("1010010001110000", '0', '1', "10", "111", "000", "100", '0', '-', "00"), -- i=6558
      ("1010110001110000", '1', '1', "10", "111", "000", "100", '0', '-', "00"), -- i=6559
      ("1010110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6560
      ("1011010001110000", '0', '1', "11", "111", "000", "100", '0', '-', "00"), -- i=6561
      ("1011110001110000", '1', '1', "11", "111", "000", "100", '0', '-', "00"), -- i=6562
      ("1011110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6563
      ("0101010001110000", '0', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6564
      ("0101110001110000", '1', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6565
      ("0101110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6566
      ("0100010001110000", '0', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6567
      ("0100110001110000", '1', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6568
      ("0100110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6569
      ("0000010000001010", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6570
      ("0000110000001010", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6571
      ("0000110000001010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6572
      ("1000010001110001", '0', '1', "00", "111", "001", "100", '0', '-', "00"), -- i=6573
      ("1000110001110001", '1', '1', "00", "111", "001", "100", '0', '-', "00"), -- i=6574
      ("1000110001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6575
      ("1001010001110001", '0', '1', "01", "111", "001", "100", '0', '-', "00"), -- i=6576
      ("1001110001110001", '1', '1', "01", "111", "001", "100", '0', '-', "00"), -- i=6577
      ("1001110001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6578
      ("1010010001110001", '0', '1', "10", "111", "001", "100", '0', '-', "00"), -- i=6579
      ("1010110001110001", '1', '1', "10", "111", "001", "100", '0', '-', "00"), -- i=6580
      ("1010110001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6581
      ("1011010001110001", '0', '1', "11", "111", "001", "100", '0', '-', "00"), -- i=6582
      ("1011110001110001", '1', '1', "11", "111", "001", "100", '0', '-', "00"), -- i=6583
      ("1011110001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6584
      ("0101010001110000", '0', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6585
      ("0101110001110000", '1', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6586
      ("0101110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6587
      ("0100010001110000", '0', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6588
      ("0100110001110000", '1', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6589
      ("0100110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6590
      ("0000010011101100", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6591
      ("0000110011101100", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6592
      ("0000110011101100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6593
      ("1000010001110010", '0', '1', "00", "111", "010", "100", '0', '-', "00"), -- i=6594
      ("1000110001110010", '1', '1', "00", "111", "010", "100", '0', '-', "00"), -- i=6595
      ("1000110001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6596
      ("1001010001110010", '0', '1', "01", "111", "010", "100", '0', '-', "00"), -- i=6597
      ("1001110001110010", '1', '1', "01", "111", "010", "100", '0', '-', "00"), -- i=6598
      ("1001110001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6599
      ("1010010001110010", '0', '1', "10", "111", "010", "100", '0', '-', "00"), -- i=6600
      ("1010110001110010", '1', '1', "10", "111", "010", "100", '0', '-', "00"), -- i=6601
      ("1010110001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6602
      ("1011010001110010", '0', '1', "11", "111", "010", "100", '0', '-', "00"), -- i=6603
      ("1011110001110010", '1', '1', "11", "111", "010", "100", '0', '-', "00"), -- i=6604
      ("1011110001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6605
      ("0101010001110000", '0', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6606
      ("0101110001110000", '1', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6607
      ("0101110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6608
      ("0100010001110000", '0', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6609
      ("0100110001110000", '1', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6610
      ("0100110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6611
      ("0000010000011100", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6612
      ("0000110000011100", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6613
      ("0000110000011100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6614
      ("1000010001110011", '0', '1', "00", "111", "011", "100", '0', '-', "00"), -- i=6615
      ("1000110001110011", '1', '1', "00", "111", "011", "100", '0', '-', "00"), -- i=6616
      ("1000110001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6617
      ("1001010001110011", '0', '1', "01", "111", "011", "100", '0', '-', "00"), -- i=6618
      ("1001110001110011", '1', '1', "01", "111", "011", "100", '0', '-', "00"), -- i=6619
      ("1001110001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6620
      ("1010010001110011", '0', '1', "10", "111", "011", "100", '0', '-', "00"), -- i=6621
      ("1010110001110011", '1', '1', "10", "111", "011", "100", '0', '-', "00"), -- i=6622
      ("1010110001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6623
      ("1011010001110011", '0', '1', "11", "111", "011", "100", '0', '-', "00"), -- i=6624
      ("1011110001110011", '1', '1', "11", "111", "011", "100", '0', '-', "00"), -- i=6625
      ("1011110001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6626
      ("0101010001110000", '0', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6627
      ("0101110001110000", '1', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6628
      ("0101110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6629
      ("0100010001110000", '0', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6630
      ("0100110001110000", '1', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6631
      ("0100110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6632
      ("0000010001000010", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6633
      ("0000110001000010", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6634
      ("0000110001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6635
      ("1000010001110100", '0', '1', "00", "111", "100", "100", '0', '-', "00"), -- i=6636
      ("1000110001110100", '1', '1', "00", "111", "100", "100", '0', '-', "00"), -- i=6637
      ("1000110001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6638
      ("1001010001110100", '0', '1', "01", "111", "100", "100", '0', '-', "00"), -- i=6639
      ("1001110001110100", '1', '1', "01", "111", "100", "100", '0', '-', "00"), -- i=6640
      ("1001110001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6641
      ("1010010001110100", '0', '1', "10", "111", "100", "100", '0', '-', "00"), -- i=6642
      ("1010110001110100", '1', '1', "10", "111", "100", "100", '0', '-', "00"), -- i=6643
      ("1010110001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6644
      ("1011010001110100", '0', '1', "11", "111", "100", "100", '0', '-', "00"), -- i=6645
      ("1011110001110100", '1', '1', "11", "111", "100", "100", '0', '-', "00"), -- i=6646
      ("1011110001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6647
      ("0101010001110000", '0', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6648
      ("0101110001110000", '1', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6649
      ("0101110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6650
      ("0100010001110000", '0', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6651
      ("0100110001110000", '1', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6652
      ("0100110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6653
      ("0000010011101101", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6654
      ("0000110011101101", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6655
      ("0000110011101101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6656
      ("1000010001110101", '0', '1', "00", "111", "101", "100", '0', '-', "00"), -- i=6657
      ("1000110001110101", '1', '1', "00", "111", "101", "100", '0', '-', "00"), -- i=6658
      ("1000110001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6659
      ("1001010001110101", '0', '1', "01", "111", "101", "100", '0', '-', "00"), -- i=6660
      ("1001110001110101", '1', '1', "01", "111", "101", "100", '0', '-', "00"), -- i=6661
      ("1001110001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6662
      ("1010010001110101", '0', '1', "10", "111", "101", "100", '0', '-', "00"), -- i=6663
      ("1010110001110101", '1', '1', "10", "111", "101", "100", '0', '-', "00"), -- i=6664
      ("1010110001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6665
      ("1011010001110101", '0', '1', "11", "111", "101", "100", '0', '-', "00"), -- i=6666
      ("1011110001110101", '1', '1', "11", "111", "101", "100", '0', '-', "00"), -- i=6667
      ("1011110001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6668
      ("0101010001110000", '0', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6669
      ("0101110001110000", '1', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6670
      ("0101110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6671
      ("0100010001110000", '0', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6672
      ("0100110001110000", '1', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6673
      ("0100110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6674
      ("0000010000000001", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6675
      ("0000110000000001", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6676
      ("0000110000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6677
      ("1000010001110110", '0', '1', "00", "111", "110", "100", '0', '-', "00"), -- i=6678
      ("1000110001110110", '1', '1', "00", "111", "110", "100", '0', '-', "00"), -- i=6679
      ("1000110001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6680
      ("1001010001110110", '0', '1', "01", "111", "110", "100", '0', '-', "00"), -- i=6681
      ("1001110001110110", '1', '1', "01", "111", "110", "100", '0', '-', "00"), -- i=6682
      ("1001110001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6683
      ("1010010001110110", '0', '1', "10", "111", "110", "100", '0', '-', "00"), -- i=6684
      ("1010110001110110", '1', '1', "10", "111", "110", "100", '0', '-', "00"), -- i=6685
      ("1010110001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6686
      ("1011010001110110", '0', '1', "11", "111", "110", "100", '0', '-', "00"), -- i=6687
      ("1011110001110110", '1', '1', "11", "111", "110", "100", '0', '-', "00"), -- i=6688
      ("1011110001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6689
      ("0101010001110000", '0', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6690
      ("0101110001110000", '1', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6691
      ("0101110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6692
      ("0100010001110000", '0', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6693
      ("0100110001110000", '1', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6694
      ("0100110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6695
      ("0000010001100111", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6696
      ("0000110001100111", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6697
      ("0000110001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6698
      ("1000010001110111", '0', '1', "00", "111", "111", "100", '0', '-', "00"), -- i=6699
      ("1000110001110111", '1', '1', "00", "111", "111", "100", '0', '-', "00"), -- i=6700
      ("1000110001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6701
      ("1001010001110111", '0', '1', "01", "111", "111", "100", '0', '-', "00"), -- i=6702
      ("1001110001110111", '1', '1', "01", "111", "111", "100", '0', '-', "00"), -- i=6703
      ("1001110001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6704
      ("1010010001110111", '0', '1', "10", "111", "111", "100", '0', '-', "00"), -- i=6705
      ("1010110001110111", '1', '1', "10", "111", "111", "100", '0', '-', "00"), -- i=6706
      ("1010110001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6707
      ("1011010001110111", '0', '1', "11", "111", "111", "100", '0', '-', "00"), -- i=6708
      ("1011110001110111", '1', '1', "11", "111", "111", "100", '0', '-', "00"), -- i=6709
      ("1011110001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6710
      ("0101010001110000", '0', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6711
      ("0101110001110000", '1', '1', "--", "111", "---", "100", '0', '1', "01"), -- i=6712
      ("0101110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6713
      ("0100010001110000", '0', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6714
      ("0100110001110000", '1', '0', "--", "111", "100", "---", '1', '-', "--"), -- i=6715
      ("0100110001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6716
      ("0000010000001110", '0', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6717
      ("0000110000001110", '1', '1', "--", "---", "---", "100", '0', '-', "10"), -- i=6718
      ("0000110000001110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6719
      ("1000010100000000", '0', '1', "00", "000", "000", "101", '0', '-', "00"), -- i=6720
      ("1000110100000000", '1', '1', "00", "000", "000", "101", '0', '-', "00"), -- i=6721
      ("1000110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6722
      ("1001010100000000", '0', '1', "01", "000", "000", "101", '0', '-', "00"), -- i=6723
      ("1001110100000000", '1', '1', "01", "000", "000", "101", '0', '-', "00"), -- i=6724
      ("1001110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6725
      ("1010010100000000", '0', '1', "10", "000", "000", "101", '0', '-', "00"), -- i=6726
      ("1010110100000000", '1', '1', "10", "000", "000", "101", '0', '-', "00"), -- i=6727
      ("1010110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6728
      ("1011010100000000", '0', '1', "11", "000", "000", "101", '0', '-', "00"), -- i=6729
      ("1011110100000000", '1', '1', "11", "000", "000", "101", '0', '-', "00"), -- i=6730
      ("1011110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6731
      ("0101010100000000", '0', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6732
      ("0101110100000000", '1', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6733
      ("0101110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6734
      ("0100010100000000", '0', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6735
      ("0100110100000000", '1', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6736
      ("0100110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6737
      ("0000010111100100", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6738
      ("0000110111100100", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6739
      ("0000110111100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6740
      ("1000010100000001", '0', '1', "00", "000", "001", "101", '0', '-', "00"), -- i=6741
      ("1000110100000001", '1', '1', "00", "000", "001", "101", '0', '-', "00"), -- i=6742
      ("1000110100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6743
      ("1001010100000001", '0', '1', "01", "000", "001", "101", '0', '-', "00"), -- i=6744
      ("1001110100000001", '1', '1', "01", "000", "001", "101", '0', '-', "00"), -- i=6745
      ("1001110100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6746
      ("1010010100000001", '0', '1', "10", "000", "001", "101", '0', '-', "00"), -- i=6747
      ("1010110100000001", '1', '1', "10", "000", "001", "101", '0', '-', "00"), -- i=6748
      ("1010110100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6749
      ("1011010100000001", '0', '1', "11", "000", "001", "101", '0', '-', "00"), -- i=6750
      ("1011110100000001", '1', '1', "11", "000", "001", "101", '0', '-', "00"), -- i=6751
      ("1011110100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6752
      ("0101010100000000", '0', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6753
      ("0101110100000000", '1', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6754
      ("0101110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6755
      ("0100010100000000", '0', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6756
      ("0100110100000000", '1', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6757
      ("0100110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6758
      ("0000010111101101", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6759
      ("0000110111101101", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6760
      ("0000110111101101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6761
      ("1000010100000010", '0', '1', "00", "000", "010", "101", '0', '-', "00"), -- i=6762
      ("1000110100000010", '1', '1', "00", "000", "010", "101", '0', '-', "00"), -- i=6763
      ("1000110100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6764
      ("1001010100000010", '0', '1', "01", "000", "010", "101", '0', '-', "00"), -- i=6765
      ("1001110100000010", '1', '1', "01", "000", "010", "101", '0', '-', "00"), -- i=6766
      ("1001110100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6767
      ("1010010100000010", '0', '1', "10", "000", "010", "101", '0', '-', "00"), -- i=6768
      ("1010110100000010", '1', '1', "10", "000", "010", "101", '0', '-', "00"), -- i=6769
      ("1010110100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6770
      ("1011010100000010", '0', '1', "11", "000", "010", "101", '0', '-', "00"), -- i=6771
      ("1011110100000010", '1', '1', "11", "000", "010", "101", '0', '-', "00"), -- i=6772
      ("1011110100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6773
      ("0101010100000000", '0', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6774
      ("0101110100000000", '1', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6775
      ("0101110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6776
      ("0100010100000000", '0', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6777
      ("0100110100000000", '1', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6778
      ("0100110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6779
      ("0000010101010001", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6780
      ("0000110101010001", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6781
      ("0000110101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6782
      ("1000010100000011", '0', '1', "00", "000", "011", "101", '0', '-', "00"), -- i=6783
      ("1000110100000011", '1', '1', "00", "000", "011", "101", '0', '-', "00"), -- i=6784
      ("1000110100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6785
      ("1001010100000011", '0', '1', "01", "000", "011", "101", '0', '-', "00"), -- i=6786
      ("1001110100000011", '1', '1', "01", "000", "011", "101", '0', '-', "00"), -- i=6787
      ("1001110100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6788
      ("1010010100000011", '0', '1', "10", "000", "011", "101", '0', '-', "00"), -- i=6789
      ("1010110100000011", '1', '1', "10", "000", "011", "101", '0', '-', "00"), -- i=6790
      ("1010110100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6791
      ("1011010100000011", '0', '1', "11", "000", "011", "101", '0', '-', "00"), -- i=6792
      ("1011110100000011", '1', '1', "11", "000", "011", "101", '0', '-', "00"), -- i=6793
      ("1011110100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6794
      ("0101010100000000", '0', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6795
      ("0101110100000000", '1', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6796
      ("0101110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6797
      ("0100010100000000", '0', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6798
      ("0100110100000000", '1', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6799
      ("0100110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6800
      ("0000010100011100", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6801
      ("0000110100011100", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6802
      ("0000110100011100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6803
      ("1000010100000100", '0', '1', "00", "000", "100", "101", '0', '-', "00"), -- i=6804
      ("1000110100000100", '1', '1', "00", "000", "100", "101", '0', '-', "00"), -- i=6805
      ("1000110100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6806
      ("1001010100000100", '0', '1', "01", "000", "100", "101", '0', '-', "00"), -- i=6807
      ("1001110100000100", '1', '1', "01", "000", "100", "101", '0', '-', "00"), -- i=6808
      ("1001110100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6809
      ("1010010100000100", '0', '1', "10", "000", "100", "101", '0', '-', "00"), -- i=6810
      ("1010110100000100", '1', '1', "10", "000", "100", "101", '0', '-', "00"), -- i=6811
      ("1010110100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6812
      ("1011010100000100", '0', '1', "11", "000", "100", "101", '0', '-', "00"), -- i=6813
      ("1011110100000100", '1', '1', "11", "000", "100", "101", '0', '-', "00"), -- i=6814
      ("1011110100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6815
      ("0101010100000000", '0', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6816
      ("0101110100000000", '1', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6817
      ("0101110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6818
      ("0100010100000000", '0', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6819
      ("0100110100000000", '1', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6820
      ("0100110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6821
      ("0000010100011011", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6822
      ("0000110100011011", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6823
      ("0000110100011011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6824
      ("1000010100000101", '0', '1', "00", "000", "101", "101", '0', '-', "00"), -- i=6825
      ("1000110100000101", '1', '1', "00", "000", "101", "101", '0', '-', "00"), -- i=6826
      ("1000110100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6827
      ("1001010100000101", '0', '1', "01", "000", "101", "101", '0', '-', "00"), -- i=6828
      ("1001110100000101", '1', '1', "01", "000", "101", "101", '0', '-', "00"), -- i=6829
      ("1001110100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6830
      ("1010010100000101", '0', '1', "10", "000", "101", "101", '0', '-', "00"), -- i=6831
      ("1010110100000101", '1', '1', "10", "000", "101", "101", '0', '-', "00"), -- i=6832
      ("1010110100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6833
      ("1011010100000101", '0', '1', "11", "000", "101", "101", '0', '-', "00"), -- i=6834
      ("1011110100000101", '1', '1', "11", "000", "101", "101", '0', '-', "00"), -- i=6835
      ("1011110100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6836
      ("0101010100000000", '0', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6837
      ("0101110100000000", '1', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6838
      ("0101110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6839
      ("0100010100000000", '0', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6840
      ("0100110100000000", '1', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6841
      ("0100110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6842
      ("0000010110110111", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6843
      ("0000110110110111", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6844
      ("0000110110110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6845
      ("1000010100000110", '0', '1', "00", "000", "110", "101", '0', '-', "00"), -- i=6846
      ("1000110100000110", '1', '1', "00", "000", "110", "101", '0', '-', "00"), -- i=6847
      ("1000110100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6848
      ("1001010100000110", '0', '1', "01", "000", "110", "101", '0', '-', "00"), -- i=6849
      ("1001110100000110", '1', '1', "01", "000", "110", "101", '0', '-', "00"), -- i=6850
      ("1001110100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6851
      ("1010010100000110", '0', '1', "10", "000", "110", "101", '0', '-', "00"), -- i=6852
      ("1010110100000110", '1', '1', "10", "000", "110", "101", '0', '-', "00"), -- i=6853
      ("1010110100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6854
      ("1011010100000110", '0', '1', "11", "000", "110", "101", '0', '-', "00"), -- i=6855
      ("1011110100000110", '1', '1', "11", "000", "110", "101", '0', '-', "00"), -- i=6856
      ("1011110100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6857
      ("0101010100000000", '0', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6858
      ("0101110100000000", '1', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6859
      ("0101110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6860
      ("0100010100000000", '0', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6861
      ("0100110100000000", '1', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6862
      ("0100110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6863
      ("0000010101011001", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6864
      ("0000110101011001", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6865
      ("0000110101011001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6866
      ("1000010100000111", '0', '1', "00", "000", "111", "101", '0', '-', "00"), -- i=6867
      ("1000110100000111", '1', '1', "00", "000", "111", "101", '0', '-', "00"), -- i=6868
      ("1000110100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6869
      ("1001010100000111", '0', '1', "01", "000", "111", "101", '0', '-', "00"), -- i=6870
      ("1001110100000111", '1', '1', "01", "000", "111", "101", '0', '-', "00"), -- i=6871
      ("1001110100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6872
      ("1010010100000111", '0', '1', "10", "000", "111", "101", '0', '-', "00"), -- i=6873
      ("1010110100000111", '1', '1', "10", "000", "111", "101", '0', '-', "00"), -- i=6874
      ("1010110100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6875
      ("1011010100000111", '0', '1', "11", "000", "111", "101", '0', '-', "00"), -- i=6876
      ("1011110100000111", '1', '1', "11", "000", "111", "101", '0', '-', "00"), -- i=6877
      ("1011110100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6878
      ("0101010100000000", '0', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6879
      ("0101110100000000", '1', '1', "--", "000", "---", "101", '0', '1', "01"), -- i=6880
      ("0101110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6881
      ("0100010100000000", '0', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6882
      ("0100110100000000", '1', '0', "--", "000", "101", "---", '1', '-', "--"), -- i=6883
      ("0100110100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6884
      ("0000010111101011", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6885
      ("0000110111101011", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6886
      ("0000110111101011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6887
      ("1000010100010000", '0', '1', "00", "001", "000", "101", '0', '-', "00"), -- i=6888
      ("1000110100010000", '1', '1', "00", "001", "000", "101", '0', '-', "00"), -- i=6889
      ("1000110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6890
      ("1001010100010000", '0', '1', "01", "001", "000", "101", '0', '-', "00"), -- i=6891
      ("1001110100010000", '1', '1', "01", "001", "000", "101", '0', '-', "00"), -- i=6892
      ("1001110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6893
      ("1010010100010000", '0', '1', "10", "001", "000", "101", '0', '-', "00"), -- i=6894
      ("1010110100010000", '1', '1', "10", "001", "000", "101", '0', '-', "00"), -- i=6895
      ("1010110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6896
      ("1011010100010000", '0', '1', "11", "001", "000", "101", '0', '-', "00"), -- i=6897
      ("1011110100010000", '1', '1', "11", "001", "000", "101", '0', '-', "00"), -- i=6898
      ("1011110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6899
      ("0101010100010000", '0', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=6900
      ("0101110100010000", '1', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=6901
      ("0101110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6902
      ("0100010100010000", '0', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=6903
      ("0100110100010000", '1', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=6904
      ("0100110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6905
      ("0000010111010100", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6906
      ("0000110111010100", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6907
      ("0000110111010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6908
      ("1000010100010001", '0', '1', "00", "001", "001", "101", '0', '-', "00"), -- i=6909
      ("1000110100010001", '1', '1', "00", "001", "001", "101", '0', '-', "00"), -- i=6910
      ("1000110100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6911
      ("1001010100010001", '0', '1', "01", "001", "001", "101", '0', '-', "00"), -- i=6912
      ("1001110100010001", '1', '1', "01", "001", "001", "101", '0', '-', "00"), -- i=6913
      ("1001110100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6914
      ("1010010100010001", '0', '1', "10", "001", "001", "101", '0', '-', "00"), -- i=6915
      ("1010110100010001", '1', '1', "10", "001", "001", "101", '0', '-', "00"), -- i=6916
      ("1010110100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6917
      ("1011010100010001", '0', '1', "11", "001", "001", "101", '0', '-', "00"), -- i=6918
      ("1011110100010001", '1', '1', "11", "001", "001", "101", '0', '-', "00"), -- i=6919
      ("1011110100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6920
      ("0101010100010000", '0', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=6921
      ("0101110100010000", '1', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=6922
      ("0101110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6923
      ("0100010100010000", '0', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=6924
      ("0100110100010000", '1', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=6925
      ("0100110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6926
      ("0000010100001100", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6927
      ("0000110100001100", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6928
      ("0000110100001100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6929
      ("1000010100010010", '0', '1', "00", "001", "010", "101", '0', '-', "00"), -- i=6930
      ("1000110100010010", '1', '1', "00", "001", "010", "101", '0', '-', "00"), -- i=6931
      ("1000110100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6932
      ("1001010100010010", '0', '1', "01", "001", "010", "101", '0', '-', "00"), -- i=6933
      ("1001110100010010", '1', '1', "01", "001", "010", "101", '0', '-', "00"), -- i=6934
      ("1001110100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6935
      ("1010010100010010", '0', '1', "10", "001", "010", "101", '0', '-', "00"), -- i=6936
      ("1010110100010010", '1', '1', "10", "001", "010", "101", '0', '-', "00"), -- i=6937
      ("1010110100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6938
      ("1011010100010010", '0', '1', "11", "001", "010", "101", '0', '-', "00"), -- i=6939
      ("1011110100010010", '1', '1', "11", "001", "010", "101", '0', '-', "00"), -- i=6940
      ("1011110100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6941
      ("0101010100010000", '0', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=6942
      ("0101110100010000", '1', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=6943
      ("0101110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6944
      ("0100010100010000", '0', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=6945
      ("0100110100010000", '1', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=6946
      ("0100110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6947
      ("0000010100011000", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6948
      ("0000110100011000", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6949
      ("0000110100011000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6950
      ("1000010100010011", '0', '1', "00", "001", "011", "101", '0', '-', "00"), -- i=6951
      ("1000110100010011", '1', '1', "00", "001", "011", "101", '0', '-', "00"), -- i=6952
      ("1000110100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6953
      ("1001010100010011", '0', '1', "01", "001", "011", "101", '0', '-', "00"), -- i=6954
      ("1001110100010011", '1', '1', "01", "001", "011", "101", '0', '-', "00"), -- i=6955
      ("1001110100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6956
      ("1010010100010011", '0', '1', "10", "001", "011", "101", '0', '-', "00"), -- i=6957
      ("1010110100010011", '1', '1', "10", "001", "011", "101", '0', '-', "00"), -- i=6958
      ("1010110100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6959
      ("1011010100010011", '0', '1', "11", "001", "011", "101", '0', '-', "00"), -- i=6960
      ("1011110100010011", '1', '1', "11", "001", "011", "101", '0', '-', "00"), -- i=6961
      ("1011110100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6962
      ("0101010100010000", '0', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=6963
      ("0101110100010000", '1', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=6964
      ("0101110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6965
      ("0100010100010000", '0', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=6966
      ("0100110100010000", '1', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=6967
      ("0100110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6968
      ("0000010111001011", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6969
      ("0000110111001011", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6970
      ("0000110111001011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6971
      ("1000010100010100", '0', '1', "00", "001", "100", "101", '0', '-', "00"), -- i=6972
      ("1000110100010100", '1', '1', "00", "001", "100", "101", '0', '-', "00"), -- i=6973
      ("1000110100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6974
      ("1001010100010100", '0', '1', "01", "001", "100", "101", '0', '-', "00"), -- i=6975
      ("1001110100010100", '1', '1', "01", "001", "100", "101", '0', '-', "00"), -- i=6976
      ("1001110100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6977
      ("1010010100010100", '0', '1', "10", "001", "100", "101", '0', '-', "00"), -- i=6978
      ("1010110100010100", '1', '1', "10", "001", "100", "101", '0', '-', "00"), -- i=6979
      ("1010110100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6980
      ("1011010100010100", '0', '1', "11", "001", "100", "101", '0', '-', "00"), -- i=6981
      ("1011110100010100", '1', '1', "11", "001", "100", "101", '0', '-', "00"), -- i=6982
      ("1011110100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6983
      ("0101010100010000", '0', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=6984
      ("0101110100010000", '1', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=6985
      ("0101110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6986
      ("0100010100010000", '0', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=6987
      ("0100110100010000", '1', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=6988
      ("0100110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6989
      ("0000010110111110", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6990
      ("0000110110111110", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=6991
      ("0000110110111110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6992
      ("1000010100010101", '0', '1', "00", "001", "101", "101", '0', '-', "00"), -- i=6993
      ("1000110100010101", '1', '1', "00", "001", "101", "101", '0', '-', "00"), -- i=6994
      ("1000110100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6995
      ("1001010100010101", '0', '1', "01", "001", "101", "101", '0', '-', "00"), -- i=6996
      ("1001110100010101", '1', '1', "01", "001", "101", "101", '0', '-', "00"), -- i=6997
      ("1001110100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=6998
      ("1010010100010101", '0', '1', "10", "001", "101", "101", '0', '-', "00"), -- i=6999
      ("1010110100010101", '1', '1', "10", "001", "101", "101", '0', '-', "00"), -- i=7000
      ("1010110100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7001
      ("1011010100010101", '0', '1', "11", "001", "101", "101", '0', '-', "00"), -- i=7002
      ("1011110100010101", '1', '1', "11", "001", "101", "101", '0', '-', "00"), -- i=7003
      ("1011110100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7004
      ("0101010100010000", '0', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=7005
      ("0101110100010000", '1', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=7006
      ("0101110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7007
      ("0100010100010000", '0', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=7008
      ("0100110100010000", '1', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=7009
      ("0100110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7010
      ("0000010101001101", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7011
      ("0000110101001101", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7012
      ("0000110101001101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7013
      ("1000010100010110", '0', '1', "00", "001", "110", "101", '0', '-', "00"), -- i=7014
      ("1000110100010110", '1', '1', "00", "001", "110", "101", '0', '-', "00"), -- i=7015
      ("1000110100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7016
      ("1001010100010110", '0', '1', "01", "001", "110", "101", '0', '-', "00"), -- i=7017
      ("1001110100010110", '1', '1', "01", "001", "110", "101", '0', '-', "00"), -- i=7018
      ("1001110100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7019
      ("1010010100010110", '0', '1', "10", "001", "110", "101", '0', '-', "00"), -- i=7020
      ("1010110100010110", '1', '1', "10", "001", "110", "101", '0', '-', "00"), -- i=7021
      ("1010110100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7022
      ("1011010100010110", '0', '1', "11", "001", "110", "101", '0', '-', "00"), -- i=7023
      ("1011110100010110", '1', '1', "11", "001", "110", "101", '0', '-', "00"), -- i=7024
      ("1011110100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7025
      ("0101010100010000", '0', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=7026
      ("0101110100010000", '1', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=7027
      ("0101110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7028
      ("0100010100010000", '0', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=7029
      ("0100110100010000", '1', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=7030
      ("0100110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7031
      ("0000010100010011", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7032
      ("0000110100010011", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7033
      ("0000110100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7034
      ("1000010100010111", '0', '1', "00", "001", "111", "101", '0', '-', "00"), -- i=7035
      ("1000110100010111", '1', '1', "00", "001", "111", "101", '0', '-', "00"), -- i=7036
      ("1000110100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7037
      ("1001010100010111", '0', '1', "01", "001", "111", "101", '0', '-', "00"), -- i=7038
      ("1001110100010111", '1', '1', "01", "001", "111", "101", '0', '-', "00"), -- i=7039
      ("1001110100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7040
      ("1010010100010111", '0', '1', "10", "001", "111", "101", '0', '-', "00"), -- i=7041
      ("1010110100010111", '1', '1', "10", "001", "111", "101", '0', '-', "00"), -- i=7042
      ("1010110100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7043
      ("1011010100010111", '0', '1', "11", "001", "111", "101", '0', '-', "00"), -- i=7044
      ("1011110100010111", '1', '1', "11", "001", "111", "101", '0', '-', "00"), -- i=7045
      ("1011110100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7046
      ("0101010100010000", '0', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=7047
      ("0101110100010000", '1', '1', "--", "001", "---", "101", '0', '1', "01"), -- i=7048
      ("0101110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7049
      ("0100010100010000", '0', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=7050
      ("0100110100010000", '1', '0', "--", "001", "101", "---", '1', '-', "--"), -- i=7051
      ("0100110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7052
      ("0000010111001110", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7053
      ("0000110111001110", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7054
      ("0000110111001110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7055
      ("1000010100100000", '0', '1', "00", "010", "000", "101", '0', '-', "00"), -- i=7056
      ("1000110100100000", '1', '1', "00", "010", "000", "101", '0', '-', "00"), -- i=7057
      ("1000110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7058
      ("1001010100100000", '0', '1', "01", "010", "000", "101", '0', '-', "00"), -- i=7059
      ("1001110100100000", '1', '1', "01", "010", "000", "101", '0', '-', "00"), -- i=7060
      ("1001110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7061
      ("1010010100100000", '0', '1', "10", "010", "000", "101", '0', '-', "00"), -- i=7062
      ("1010110100100000", '1', '1', "10", "010", "000", "101", '0', '-', "00"), -- i=7063
      ("1010110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7064
      ("1011010100100000", '0', '1', "11", "010", "000", "101", '0', '-', "00"), -- i=7065
      ("1011110100100000", '1', '1', "11", "010", "000", "101", '0', '-', "00"), -- i=7066
      ("1011110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7067
      ("0101010100100000", '0', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7068
      ("0101110100100000", '1', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7069
      ("0101110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7070
      ("0100010100100000", '0', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7071
      ("0100110100100000", '1', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7072
      ("0100110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7073
      ("0000010110110111", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7074
      ("0000110110110111", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7075
      ("0000110110110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7076
      ("1000010100100001", '0', '1', "00", "010", "001", "101", '0', '-', "00"), -- i=7077
      ("1000110100100001", '1', '1', "00", "010", "001", "101", '0', '-', "00"), -- i=7078
      ("1000110100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7079
      ("1001010100100001", '0', '1', "01", "010", "001", "101", '0', '-', "00"), -- i=7080
      ("1001110100100001", '1', '1', "01", "010", "001", "101", '0', '-', "00"), -- i=7081
      ("1001110100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7082
      ("1010010100100001", '0', '1', "10", "010", "001", "101", '0', '-', "00"), -- i=7083
      ("1010110100100001", '1', '1', "10", "010", "001", "101", '0', '-', "00"), -- i=7084
      ("1010110100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7085
      ("1011010100100001", '0', '1', "11", "010", "001", "101", '0', '-', "00"), -- i=7086
      ("1011110100100001", '1', '1', "11", "010", "001", "101", '0', '-', "00"), -- i=7087
      ("1011110100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7088
      ("0101010100100000", '0', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7089
      ("0101110100100000", '1', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7090
      ("0101110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7091
      ("0100010100100000", '0', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7092
      ("0100110100100000", '1', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7093
      ("0100110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7094
      ("0000010110010111", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7095
      ("0000110110010111", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7096
      ("0000110110010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7097
      ("1000010100100010", '0', '1', "00", "010", "010", "101", '0', '-', "00"), -- i=7098
      ("1000110100100010", '1', '1', "00", "010", "010", "101", '0', '-', "00"), -- i=7099
      ("1000110100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7100
      ("1001010100100010", '0', '1', "01", "010", "010", "101", '0', '-', "00"), -- i=7101
      ("1001110100100010", '1', '1', "01", "010", "010", "101", '0', '-', "00"), -- i=7102
      ("1001110100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7103
      ("1010010100100010", '0', '1', "10", "010", "010", "101", '0', '-', "00"), -- i=7104
      ("1010110100100010", '1', '1', "10", "010", "010", "101", '0', '-', "00"), -- i=7105
      ("1010110100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7106
      ("1011010100100010", '0', '1', "11", "010", "010", "101", '0', '-', "00"), -- i=7107
      ("1011110100100010", '1', '1', "11", "010", "010", "101", '0', '-', "00"), -- i=7108
      ("1011110100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7109
      ("0101010100100000", '0', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7110
      ("0101110100100000", '1', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7111
      ("0101110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7112
      ("0100010100100000", '0', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7113
      ("0100110100100000", '1', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7114
      ("0100110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7115
      ("0000010111011000", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7116
      ("0000110111011000", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7117
      ("0000110111011000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7118
      ("1000010100100011", '0', '1', "00", "010", "011", "101", '0', '-', "00"), -- i=7119
      ("1000110100100011", '1', '1', "00", "010", "011", "101", '0', '-', "00"), -- i=7120
      ("1000110100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7121
      ("1001010100100011", '0', '1', "01", "010", "011", "101", '0', '-', "00"), -- i=7122
      ("1001110100100011", '1', '1', "01", "010", "011", "101", '0', '-', "00"), -- i=7123
      ("1001110100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7124
      ("1010010100100011", '0', '1', "10", "010", "011", "101", '0', '-', "00"), -- i=7125
      ("1010110100100011", '1', '1', "10", "010", "011", "101", '0', '-', "00"), -- i=7126
      ("1010110100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7127
      ("1011010100100011", '0', '1', "11", "010", "011", "101", '0', '-', "00"), -- i=7128
      ("1011110100100011", '1', '1', "11", "010", "011", "101", '0', '-', "00"), -- i=7129
      ("1011110100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7130
      ("0101010100100000", '0', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7131
      ("0101110100100000", '1', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7132
      ("0101110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7133
      ("0100010100100000", '0', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7134
      ("0100110100100000", '1', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7135
      ("0100110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7136
      ("0000010110000110", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7137
      ("0000110110000110", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7138
      ("0000110110000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7139
      ("1000010100100100", '0', '1', "00", "010", "100", "101", '0', '-', "00"), -- i=7140
      ("1000110100100100", '1', '1', "00", "010", "100", "101", '0', '-', "00"), -- i=7141
      ("1000110100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7142
      ("1001010100100100", '0', '1', "01", "010", "100", "101", '0', '-', "00"), -- i=7143
      ("1001110100100100", '1', '1', "01", "010", "100", "101", '0', '-', "00"), -- i=7144
      ("1001110100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7145
      ("1010010100100100", '0', '1', "10", "010", "100", "101", '0', '-', "00"), -- i=7146
      ("1010110100100100", '1', '1', "10", "010", "100", "101", '0', '-', "00"), -- i=7147
      ("1010110100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7148
      ("1011010100100100", '0', '1', "11", "010", "100", "101", '0', '-', "00"), -- i=7149
      ("1011110100100100", '1', '1', "11", "010", "100", "101", '0', '-', "00"), -- i=7150
      ("1011110100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7151
      ("0101010100100000", '0', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7152
      ("0101110100100000", '1', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7153
      ("0101110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7154
      ("0100010100100000", '0', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7155
      ("0100110100100000", '1', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7156
      ("0100110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7157
      ("0000010100000010", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7158
      ("0000110100000010", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7159
      ("0000110100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7160
      ("1000010100100101", '0', '1', "00", "010", "101", "101", '0', '-', "00"), -- i=7161
      ("1000110100100101", '1', '1', "00", "010", "101", "101", '0', '-', "00"), -- i=7162
      ("1000110100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7163
      ("1001010100100101", '0', '1', "01", "010", "101", "101", '0', '-', "00"), -- i=7164
      ("1001110100100101", '1', '1', "01", "010", "101", "101", '0', '-', "00"), -- i=7165
      ("1001110100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7166
      ("1010010100100101", '0', '1', "10", "010", "101", "101", '0', '-', "00"), -- i=7167
      ("1010110100100101", '1', '1', "10", "010", "101", "101", '0', '-', "00"), -- i=7168
      ("1010110100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7169
      ("1011010100100101", '0', '1', "11", "010", "101", "101", '0', '-', "00"), -- i=7170
      ("1011110100100101", '1', '1', "11", "010", "101", "101", '0', '-', "00"), -- i=7171
      ("1011110100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7172
      ("0101010100100000", '0', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7173
      ("0101110100100000", '1', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7174
      ("0101110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7175
      ("0100010100100000", '0', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7176
      ("0100110100100000", '1', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7177
      ("0100110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7178
      ("0000010110011111", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7179
      ("0000110110011111", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7180
      ("0000110110011111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7181
      ("1000010100100110", '0', '1', "00", "010", "110", "101", '0', '-', "00"), -- i=7182
      ("1000110100100110", '1', '1', "00", "010", "110", "101", '0', '-', "00"), -- i=7183
      ("1000110100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7184
      ("1001010100100110", '0', '1', "01", "010", "110", "101", '0', '-', "00"), -- i=7185
      ("1001110100100110", '1', '1', "01", "010", "110", "101", '0', '-', "00"), -- i=7186
      ("1001110100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7187
      ("1010010100100110", '0', '1', "10", "010", "110", "101", '0', '-', "00"), -- i=7188
      ("1010110100100110", '1', '1', "10", "010", "110", "101", '0', '-', "00"), -- i=7189
      ("1010110100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7190
      ("1011010100100110", '0', '1', "11", "010", "110", "101", '0', '-', "00"), -- i=7191
      ("1011110100100110", '1', '1', "11", "010", "110", "101", '0', '-', "00"), -- i=7192
      ("1011110100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7193
      ("0101010100100000", '0', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7194
      ("0101110100100000", '1', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7195
      ("0101110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7196
      ("0100010100100000", '0', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7197
      ("0100110100100000", '1', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7198
      ("0100110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7199
      ("0000010101011011", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7200
      ("0000110101011011", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7201
      ("0000110101011011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7202
      ("1000010100100111", '0', '1', "00", "010", "111", "101", '0', '-', "00"), -- i=7203
      ("1000110100100111", '1', '1', "00", "010", "111", "101", '0', '-', "00"), -- i=7204
      ("1000110100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7205
      ("1001010100100111", '0', '1', "01", "010", "111", "101", '0', '-', "00"), -- i=7206
      ("1001110100100111", '1', '1', "01", "010", "111", "101", '0', '-', "00"), -- i=7207
      ("1001110100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7208
      ("1010010100100111", '0', '1', "10", "010", "111", "101", '0', '-', "00"), -- i=7209
      ("1010110100100111", '1', '1', "10", "010", "111", "101", '0', '-', "00"), -- i=7210
      ("1010110100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7211
      ("1011010100100111", '0', '1', "11", "010", "111", "101", '0', '-', "00"), -- i=7212
      ("1011110100100111", '1', '1', "11", "010", "111", "101", '0', '-', "00"), -- i=7213
      ("1011110100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7214
      ("0101010100100000", '0', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7215
      ("0101110100100000", '1', '1', "--", "010", "---", "101", '0', '1', "01"), -- i=7216
      ("0101110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7217
      ("0100010100100000", '0', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7218
      ("0100110100100000", '1', '0', "--", "010", "101", "---", '1', '-', "--"), -- i=7219
      ("0100110100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7220
      ("0000010110101110", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7221
      ("0000110110101110", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7222
      ("0000110110101110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7223
      ("1000010100110000", '0', '1', "00", "011", "000", "101", '0', '-', "00"), -- i=7224
      ("1000110100110000", '1', '1', "00", "011", "000", "101", '0', '-', "00"), -- i=7225
      ("1000110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7226
      ("1001010100110000", '0', '1', "01", "011", "000", "101", '0', '-', "00"), -- i=7227
      ("1001110100110000", '1', '1', "01", "011", "000", "101", '0', '-', "00"), -- i=7228
      ("1001110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7229
      ("1010010100110000", '0', '1', "10", "011", "000", "101", '0', '-', "00"), -- i=7230
      ("1010110100110000", '1', '1', "10", "011", "000", "101", '0', '-', "00"), -- i=7231
      ("1010110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7232
      ("1011010100110000", '0', '1', "11", "011", "000", "101", '0', '-', "00"), -- i=7233
      ("1011110100110000", '1', '1', "11", "011", "000", "101", '0', '-', "00"), -- i=7234
      ("1011110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7235
      ("0101010100110000", '0', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7236
      ("0101110100110000", '1', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7237
      ("0101110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7238
      ("0100010100110000", '0', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7239
      ("0100110100110000", '1', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7240
      ("0100110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7241
      ("0000010101000100", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7242
      ("0000110101000100", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7243
      ("0000110101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7244
      ("1000010100110001", '0', '1', "00", "011", "001", "101", '0', '-', "00"), -- i=7245
      ("1000110100110001", '1', '1', "00", "011", "001", "101", '0', '-', "00"), -- i=7246
      ("1000110100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7247
      ("1001010100110001", '0', '1', "01", "011", "001", "101", '0', '-', "00"), -- i=7248
      ("1001110100110001", '1', '1', "01", "011", "001", "101", '0', '-', "00"), -- i=7249
      ("1001110100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7250
      ("1010010100110001", '0', '1', "10", "011", "001", "101", '0', '-', "00"), -- i=7251
      ("1010110100110001", '1', '1', "10", "011", "001", "101", '0', '-', "00"), -- i=7252
      ("1010110100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7253
      ("1011010100110001", '0', '1', "11", "011", "001", "101", '0', '-', "00"), -- i=7254
      ("1011110100110001", '1', '1', "11", "011", "001", "101", '0', '-', "00"), -- i=7255
      ("1011110100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7256
      ("0101010100110000", '0', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7257
      ("0101110100110000", '1', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7258
      ("0101110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7259
      ("0100010100110000", '0', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7260
      ("0100110100110000", '1', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7261
      ("0100110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7262
      ("0000010101011110", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7263
      ("0000110101011110", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7264
      ("0000110101011110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7265
      ("1000010100110010", '0', '1', "00", "011", "010", "101", '0', '-', "00"), -- i=7266
      ("1000110100110010", '1', '1', "00", "011", "010", "101", '0', '-', "00"), -- i=7267
      ("1000110100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7268
      ("1001010100110010", '0', '1', "01", "011", "010", "101", '0', '-', "00"), -- i=7269
      ("1001110100110010", '1', '1', "01", "011", "010", "101", '0', '-', "00"), -- i=7270
      ("1001110100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7271
      ("1010010100110010", '0', '1', "10", "011", "010", "101", '0', '-', "00"), -- i=7272
      ("1010110100110010", '1', '1', "10", "011", "010", "101", '0', '-', "00"), -- i=7273
      ("1010110100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7274
      ("1011010100110010", '0', '1', "11", "011", "010", "101", '0', '-', "00"), -- i=7275
      ("1011110100110010", '1', '1', "11", "011", "010", "101", '0', '-', "00"), -- i=7276
      ("1011110100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7277
      ("0101010100110000", '0', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7278
      ("0101110100110000", '1', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7279
      ("0101110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7280
      ("0100010100110000", '0', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7281
      ("0100110100110000", '1', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7282
      ("0100110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7283
      ("0000010110100011", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7284
      ("0000110110100011", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7285
      ("0000110110100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7286
      ("1000010100110011", '0', '1', "00", "011", "011", "101", '0', '-', "00"), -- i=7287
      ("1000110100110011", '1', '1', "00", "011", "011", "101", '0', '-', "00"), -- i=7288
      ("1000110100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7289
      ("1001010100110011", '0', '1', "01", "011", "011", "101", '0', '-', "00"), -- i=7290
      ("1001110100110011", '1', '1', "01", "011", "011", "101", '0', '-', "00"), -- i=7291
      ("1001110100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7292
      ("1010010100110011", '0', '1', "10", "011", "011", "101", '0', '-', "00"), -- i=7293
      ("1010110100110011", '1', '1', "10", "011", "011", "101", '0', '-', "00"), -- i=7294
      ("1010110100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7295
      ("1011010100110011", '0', '1', "11", "011", "011", "101", '0', '-', "00"), -- i=7296
      ("1011110100110011", '1', '1', "11", "011", "011", "101", '0', '-', "00"), -- i=7297
      ("1011110100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7298
      ("0101010100110000", '0', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7299
      ("0101110100110000", '1', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7300
      ("0101110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7301
      ("0100010100110000", '0', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7302
      ("0100110100110000", '1', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7303
      ("0100110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7304
      ("0000010110111000", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7305
      ("0000110110111000", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7306
      ("0000110110111000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7307
      ("1000010100110100", '0', '1', "00", "011", "100", "101", '0', '-', "00"), -- i=7308
      ("1000110100110100", '1', '1', "00", "011", "100", "101", '0', '-', "00"), -- i=7309
      ("1000110100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7310
      ("1001010100110100", '0', '1', "01", "011", "100", "101", '0', '-', "00"), -- i=7311
      ("1001110100110100", '1', '1', "01", "011", "100", "101", '0', '-', "00"), -- i=7312
      ("1001110100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7313
      ("1010010100110100", '0', '1', "10", "011", "100", "101", '0', '-', "00"), -- i=7314
      ("1010110100110100", '1', '1', "10", "011", "100", "101", '0', '-', "00"), -- i=7315
      ("1010110100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7316
      ("1011010100110100", '0', '1', "11", "011", "100", "101", '0', '-', "00"), -- i=7317
      ("1011110100110100", '1', '1', "11", "011", "100", "101", '0', '-', "00"), -- i=7318
      ("1011110100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7319
      ("0101010100110000", '0', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7320
      ("0101110100110000", '1', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7321
      ("0101110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7322
      ("0100010100110000", '0', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7323
      ("0100110100110000", '1', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7324
      ("0100110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7325
      ("0000010111101110", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7326
      ("0000110111101110", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7327
      ("0000110111101110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7328
      ("1000010100110101", '0', '1', "00", "011", "101", "101", '0', '-', "00"), -- i=7329
      ("1000110100110101", '1', '1', "00", "011", "101", "101", '0', '-', "00"), -- i=7330
      ("1000110100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7331
      ("1001010100110101", '0', '1', "01", "011", "101", "101", '0', '-', "00"), -- i=7332
      ("1001110100110101", '1', '1', "01", "011", "101", "101", '0', '-', "00"), -- i=7333
      ("1001110100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7334
      ("1010010100110101", '0', '1', "10", "011", "101", "101", '0', '-', "00"), -- i=7335
      ("1010110100110101", '1', '1', "10", "011", "101", "101", '0', '-', "00"), -- i=7336
      ("1010110100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7337
      ("1011010100110101", '0', '1', "11", "011", "101", "101", '0', '-', "00"), -- i=7338
      ("1011110100110101", '1', '1', "11", "011", "101", "101", '0', '-', "00"), -- i=7339
      ("1011110100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7340
      ("0101010100110000", '0', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7341
      ("0101110100110000", '1', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7342
      ("0101110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7343
      ("0100010100110000", '0', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7344
      ("0100110100110000", '1', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7345
      ("0100110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7346
      ("0000010110100000", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7347
      ("0000110110100000", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7348
      ("0000110110100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7349
      ("1000010100110110", '0', '1', "00", "011", "110", "101", '0', '-', "00"), -- i=7350
      ("1000110100110110", '1', '1', "00", "011", "110", "101", '0', '-', "00"), -- i=7351
      ("1000110100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7352
      ("1001010100110110", '0', '1', "01", "011", "110", "101", '0', '-', "00"), -- i=7353
      ("1001110100110110", '1', '1', "01", "011", "110", "101", '0', '-', "00"), -- i=7354
      ("1001110100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7355
      ("1010010100110110", '0', '1', "10", "011", "110", "101", '0', '-', "00"), -- i=7356
      ("1010110100110110", '1', '1', "10", "011", "110", "101", '0', '-', "00"), -- i=7357
      ("1010110100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7358
      ("1011010100110110", '0', '1', "11", "011", "110", "101", '0', '-', "00"), -- i=7359
      ("1011110100110110", '1', '1', "11", "011", "110", "101", '0', '-', "00"), -- i=7360
      ("1011110100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7361
      ("0101010100110000", '0', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7362
      ("0101110100110000", '1', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7363
      ("0101110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7364
      ("0100010100110000", '0', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7365
      ("0100110100110000", '1', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7366
      ("0100110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7367
      ("0000010111101100", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7368
      ("0000110111101100", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7369
      ("0000110111101100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7370
      ("1000010100110111", '0', '1', "00", "011", "111", "101", '0', '-', "00"), -- i=7371
      ("1000110100110111", '1', '1', "00", "011", "111", "101", '0', '-', "00"), -- i=7372
      ("1000110100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7373
      ("1001010100110111", '0', '1', "01", "011", "111", "101", '0', '-', "00"), -- i=7374
      ("1001110100110111", '1', '1', "01", "011", "111", "101", '0', '-', "00"), -- i=7375
      ("1001110100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7376
      ("1010010100110111", '0', '1', "10", "011", "111", "101", '0', '-', "00"), -- i=7377
      ("1010110100110111", '1', '1', "10", "011", "111", "101", '0', '-', "00"), -- i=7378
      ("1010110100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7379
      ("1011010100110111", '0', '1', "11", "011", "111", "101", '0', '-', "00"), -- i=7380
      ("1011110100110111", '1', '1', "11", "011", "111", "101", '0', '-', "00"), -- i=7381
      ("1011110100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7382
      ("0101010100110000", '0', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7383
      ("0101110100110000", '1', '1', "--", "011", "---", "101", '0', '1', "01"), -- i=7384
      ("0101110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7385
      ("0100010100110000", '0', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7386
      ("0100110100110000", '1', '0', "--", "011", "101", "---", '1', '-', "--"), -- i=7387
      ("0100110100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7388
      ("0000010101100100", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7389
      ("0000110101100100", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7390
      ("0000110101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7391
      ("1000010101000000", '0', '1', "00", "100", "000", "101", '0', '-', "00"), -- i=7392
      ("1000110101000000", '1', '1', "00", "100", "000", "101", '0', '-', "00"), -- i=7393
      ("1000110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7394
      ("1001010101000000", '0', '1', "01", "100", "000", "101", '0', '-', "00"), -- i=7395
      ("1001110101000000", '1', '1', "01", "100", "000", "101", '0', '-', "00"), -- i=7396
      ("1001110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7397
      ("1010010101000000", '0', '1', "10", "100", "000", "101", '0', '-', "00"), -- i=7398
      ("1010110101000000", '1', '1', "10", "100", "000", "101", '0', '-', "00"), -- i=7399
      ("1010110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7400
      ("1011010101000000", '0', '1', "11", "100", "000", "101", '0', '-', "00"), -- i=7401
      ("1011110101000000", '1', '1', "11", "100", "000", "101", '0', '-', "00"), -- i=7402
      ("1011110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7403
      ("0101010101000000", '0', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7404
      ("0101110101000000", '1', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7405
      ("0101110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7406
      ("0100010101000000", '0', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7407
      ("0100110101000000", '1', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7408
      ("0100110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7409
      ("0000010101110011", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7410
      ("0000110101110011", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7411
      ("0000110101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7412
      ("1000010101000001", '0', '1', "00", "100", "001", "101", '0', '-', "00"), -- i=7413
      ("1000110101000001", '1', '1', "00", "100", "001", "101", '0', '-', "00"), -- i=7414
      ("1000110101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7415
      ("1001010101000001", '0', '1', "01", "100", "001", "101", '0', '-', "00"), -- i=7416
      ("1001110101000001", '1', '1', "01", "100", "001", "101", '0', '-', "00"), -- i=7417
      ("1001110101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7418
      ("1010010101000001", '0', '1', "10", "100", "001", "101", '0', '-', "00"), -- i=7419
      ("1010110101000001", '1', '1', "10", "100", "001", "101", '0', '-', "00"), -- i=7420
      ("1010110101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7421
      ("1011010101000001", '0', '1', "11", "100", "001", "101", '0', '-', "00"), -- i=7422
      ("1011110101000001", '1', '1', "11", "100", "001", "101", '0', '-', "00"), -- i=7423
      ("1011110101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7424
      ("0101010101000000", '0', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7425
      ("0101110101000000", '1', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7426
      ("0101110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7427
      ("0100010101000000", '0', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7428
      ("0100110101000000", '1', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7429
      ("0100110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7430
      ("0000010111001110", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7431
      ("0000110111001110", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7432
      ("0000110111001110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7433
      ("1000010101000010", '0', '1', "00", "100", "010", "101", '0', '-', "00"), -- i=7434
      ("1000110101000010", '1', '1', "00", "100", "010", "101", '0', '-', "00"), -- i=7435
      ("1000110101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7436
      ("1001010101000010", '0', '1', "01", "100", "010", "101", '0', '-', "00"), -- i=7437
      ("1001110101000010", '1', '1', "01", "100", "010", "101", '0', '-', "00"), -- i=7438
      ("1001110101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7439
      ("1010010101000010", '0', '1', "10", "100", "010", "101", '0', '-', "00"), -- i=7440
      ("1010110101000010", '1', '1', "10", "100", "010", "101", '0', '-', "00"), -- i=7441
      ("1010110101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7442
      ("1011010101000010", '0', '1', "11", "100", "010", "101", '0', '-', "00"), -- i=7443
      ("1011110101000010", '1', '1', "11", "100", "010", "101", '0', '-', "00"), -- i=7444
      ("1011110101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7445
      ("0101010101000000", '0', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7446
      ("0101110101000000", '1', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7447
      ("0101110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7448
      ("0100010101000000", '0', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7449
      ("0100110101000000", '1', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7450
      ("0100110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7451
      ("0000010111110010", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7452
      ("0000110111110010", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7453
      ("0000110111110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7454
      ("1000010101000011", '0', '1', "00", "100", "011", "101", '0', '-', "00"), -- i=7455
      ("1000110101000011", '1', '1', "00", "100", "011", "101", '0', '-', "00"), -- i=7456
      ("1000110101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7457
      ("1001010101000011", '0', '1', "01", "100", "011", "101", '0', '-', "00"), -- i=7458
      ("1001110101000011", '1', '1', "01", "100", "011", "101", '0', '-', "00"), -- i=7459
      ("1001110101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7460
      ("1010010101000011", '0', '1', "10", "100", "011", "101", '0', '-', "00"), -- i=7461
      ("1010110101000011", '1', '1', "10", "100", "011", "101", '0', '-', "00"), -- i=7462
      ("1010110101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7463
      ("1011010101000011", '0', '1', "11", "100", "011", "101", '0', '-', "00"), -- i=7464
      ("1011110101000011", '1', '1', "11", "100", "011", "101", '0', '-', "00"), -- i=7465
      ("1011110101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7466
      ("0101010101000000", '0', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7467
      ("0101110101000000", '1', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7468
      ("0101110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7469
      ("0100010101000000", '0', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7470
      ("0100110101000000", '1', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7471
      ("0100110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7472
      ("0000010101101011", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7473
      ("0000110101101011", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7474
      ("0000110101101011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7475
      ("1000010101000100", '0', '1', "00", "100", "100", "101", '0', '-', "00"), -- i=7476
      ("1000110101000100", '1', '1', "00", "100", "100", "101", '0', '-', "00"), -- i=7477
      ("1000110101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7478
      ("1001010101000100", '0', '1', "01", "100", "100", "101", '0', '-', "00"), -- i=7479
      ("1001110101000100", '1', '1', "01", "100", "100", "101", '0', '-', "00"), -- i=7480
      ("1001110101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7481
      ("1010010101000100", '0', '1', "10", "100", "100", "101", '0', '-', "00"), -- i=7482
      ("1010110101000100", '1', '1', "10", "100", "100", "101", '0', '-', "00"), -- i=7483
      ("1010110101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7484
      ("1011010101000100", '0', '1', "11", "100", "100", "101", '0', '-', "00"), -- i=7485
      ("1011110101000100", '1', '1', "11", "100", "100", "101", '0', '-', "00"), -- i=7486
      ("1011110101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7487
      ("0101010101000000", '0', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7488
      ("0101110101000000", '1', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7489
      ("0101110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7490
      ("0100010101000000", '0', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7491
      ("0100110101000000", '1', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7492
      ("0100110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7493
      ("0000010110101010", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7494
      ("0000110110101010", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7495
      ("0000110110101010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7496
      ("1000010101000101", '0', '1', "00", "100", "101", "101", '0', '-', "00"), -- i=7497
      ("1000110101000101", '1', '1', "00", "100", "101", "101", '0', '-', "00"), -- i=7498
      ("1000110101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7499
      ("1001010101000101", '0', '1', "01", "100", "101", "101", '0', '-', "00"), -- i=7500
      ("1001110101000101", '1', '1', "01", "100", "101", "101", '0', '-', "00"), -- i=7501
      ("1001110101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7502
      ("1010010101000101", '0', '1', "10", "100", "101", "101", '0', '-', "00"), -- i=7503
      ("1010110101000101", '1', '1', "10", "100", "101", "101", '0', '-', "00"), -- i=7504
      ("1010110101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7505
      ("1011010101000101", '0', '1', "11", "100", "101", "101", '0', '-', "00"), -- i=7506
      ("1011110101000101", '1', '1', "11", "100", "101", "101", '0', '-', "00"), -- i=7507
      ("1011110101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7508
      ("0101010101000000", '0', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7509
      ("0101110101000000", '1', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7510
      ("0101110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7511
      ("0100010101000000", '0', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7512
      ("0100110101000000", '1', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7513
      ("0100110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7514
      ("0000010101101000", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7515
      ("0000110101101000", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7516
      ("0000110101101000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7517
      ("1000010101000110", '0', '1', "00", "100", "110", "101", '0', '-', "00"), -- i=7518
      ("1000110101000110", '1', '1', "00", "100", "110", "101", '0', '-', "00"), -- i=7519
      ("1000110101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7520
      ("1001010101000110", '0', '1', "01", "100", "110", "101", '0', '-', "00"), -- i=7521
      ("1001110101000110", '1', '1', "01", "100", "110", "101", '0', '-', "00"), -- i=7522
      ("1001110101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7523
      ("1010010101000110", '0', '1', "10", "100", "110", "101", '0', '-', "00"), -- i=7524
      ("1010110101000110", '1', '1', "10", "100", "110", "101", '0', '-', "00"), -- i=7525
      ("1010110101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7526
      ("1011010101000110", '0', '1', "11", "100", "110", "101", '0', '-', "00"), -- i=7527
      ("1011110101000110", '1', '1', "11", "100", "110", "101", '0', '-', "00"), -- i=7528
      ("1011110101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7529
      ("0101010101000000", '0', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7530
      ("0101110101000000", '1', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7531
      ("0101110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7532
      ("0100010101000000", '0', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7533
      ("0100110101000000", '1', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7534
      ("0100110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7535
      ("0000010110101111", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7536
      ("0000110110101111", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7537
      ("0000110110101111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7538
      ("1000010101000111", '0', '1', "00", "100", "111", "101", '0', '-', "00"), -- i=7539
      ("1000110101000111", '1', '1', "00", "100", "111", "101", '0', '-', "00"), -- i=7540
      ("1000110101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7541
      ("1001010101000111", '0', '1', "01", "100", "111", "101", '0', '-', "00"), -- i=7542
      ("1001110101000111", '1', '1', "01", "100", "111", "101", '0', '-', "00"), -- i=7543
      ("1001110101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7544
      ("1010010101000111", '0', '1', "10", "100", "111", "101", '0', '-', "00"), -- i=7545
      ("1010110101000111", '1', '1', "10", "100", "111", "101", '0', '-', "00"), -- i=7546
      ("1010110101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7547
      ("1011010101000111", '0', '1', "11", "100", "111", "101", '0', '-', "00"), -- i=7548
      ("1011110101000111", '1', '1', "11", "100", "111", "101", '0', '-', "00"), -- i=7549
      ("1011110101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7550
      ("0101010101000000", '0', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7551
      ("0101110101000000", '1', '1', "--", "100", "---", "101", '0', '1', "01"), -- i=7552
      ("0101110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7553
      ("0100010101000000", '0', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7554
      ("0100110101000000", '1', '0', "--", "100", "101", "---", '1', '-', "--"), -- i=7555
      ("0100110101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7556
      ("0000010110011110", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7557
      ("0000110110011110", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7558
      ("0000110110011110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7559
      ("1000010101010000", '0', '1', "00", "101", "000", "101", '0', '-', "00"), -- i=7560
      ("1000110101010000", '1', '1', "00", "101", "000", "101", '0', '-', "00"), -- i=7561
      ("1000110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7562
      ("1001010101010000", '0', '1', "01", "101", "000", "101", '0', '-', "00"), -- i=7563
      ("1001110101010000", '1', '1', "01", "101", "000", "101", '0', '-', "00"), -- i=7564
      ("1001110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7565
      ("1010010101010000", '0', '1', "10", "101", "000", "101", '0', '-', "00"), -- i=7566
      ("1010110101010000", '1', '1', "10", "101", "000", "101", '0', '-', "00"), -- i=7567
      ("1010110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7568
      ("1011010101010000", '0', '1', "11", "101", "000", "101", '0', '-', "00"), -- i=7569
      ("1011110101010000", '1', '1', "11", "101", "000", "101", '0', '-', "00"), -- i=7570
      ("1011110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7571
      ("0101010101010000", '0', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7572
      ("0101110101010000", '1', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7573
      ("0101110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7574
      ("0100010101010000", '0', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7575
      ("0100110101010000", '1', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7576
      ("0100110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7577
      ("0000010111111110", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7578
      ("0000110111111110", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7579
      ("0000110111111110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7580
      ("1000010101010001", '0', '1', "00", "101", "001", "101", '0', '-', "00"), -- i=7581
      ("1000110101010001", '1', '1', "00", "101", "001", "101", '0', '-', "00"), -- i=7582
      ("1000110101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7583
      ("1001010101010001", '0', '1', "01", "101", "001", "101", '0', '-', "00"), -- i=7584
      ("1001110101010001", '1', '1', "01", "101", "001", "101", '0', '-', "00"), -- i=7585
      ("1001110101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7586
      ("1010010101010001", '0', '1', "10", "101", "001", "101", '0', '-', "00"), -- i=7587
      ("1010110101010001", '1', '1', "10", "101", "001", "101", '0', '-', "00"), -- i=7588
      ("1010110101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7589
      ("1011010101010001", '0', '1', "11", "101", "001", "101", '0', '-', "00"), -- i=7590
      ("1011110101010001", '1', '1', "11", "101", "001", "101", '0', '-', "00"), -- i=7591
      ("1011110101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7592
      ("0101010101010000", '0', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7593
      ("0101110101010000", '1', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7594
      ("0101110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7595
      ("0100010101010000", '0', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7596
      ("0100110101010000", '1', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7597
      ("0100110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7598
      ("0000010111111101", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7599
      ("0000110111111101", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7600
      ("0000110111111101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7601
      ("1000010101010010", '0', '1', "00", "101", "010", "101", '0', '-', "00"), -- i=7602
      ("1000110101010010", '1', '1', "00", "101", "010", "101", '0', '-', "00"), -- i=7603
      ("1000110101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7604
      ("1001010101010010", '0', '1', "01", "101", "010", "101", '0', '-', "00"), -- i=7605
      ("1001110101010010", '1', '1', "01", "101", "010", "101", '0', '-', "00"), -- i=7606
      ("1001110101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7607
      ("1010010101010010", '0', '1', "10", "101", "010", "101", '0', '-', "00"), -- i=7608
      ("1010110101010010", '1', '1', "10", "101", "010", "101", '0', '-', "00"), -- i=7609
      ("1010110101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7610
      ("1011010101010010", '0', '1', "11", "101", "010", "101", '0', '-', "00"), -- i=7611
      ("1011110101010010", '1', '1', "11", "101", "010", "101", '0', '-', "00"), -- i=7612
      ("1011110101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7613
      ("0101010101010000", '0', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7614
      ("0101110101010000", '1', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7615
      ("0101110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7616
      ("0100010101010000", '0', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7617
      ("0100110101010000", '1', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7618
      ("0100110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7619
      ("0000010100100101", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7620
      ("0000110100100101", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7621
      ("0000110100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7622
      ("1000010101010011", '0', '1', "00", "101", "011", "101", '0', '-', "00"), -- i=7623
      ("1000110101010011", '1', '1', "00", "101", "011", "101", '0', '-', "00"), -- i=7624
      ("1000110101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7625
      ("1001010101010011", '0', '1', "01", "101", "011", "101", '0', '-', "00"), -- i=7626
      ("1001110101010011", '1', '1', "01", "101", "011", "101", '0', '-', "00"), -- i=7627
      ("1001110101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7628
      ("1010010101010011", '0', '1', "10", "101", "011", "101", '0', '-', "00"), -- i=7629
      ("1010110101010011", '1', '1', "10", "101", "011", "101", '0', '-', "00"), -- i=7630
      ("1010110101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7631
      ("1011010101010011", '0', '1', "11", "101", "011", "101", '0', '-', "00"), -- i=7632
      ("1011110101010011", '1', '1', "11", "101", "011", "101", '0', '-', "00"), -- i=7633
      ("1011110101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7634
      ("0101010101010000", '0', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7635
      ("0101110101010000", '1', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7636
      ("0101110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7637
      ("0100010101010000", '0', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7638
      ("0100110101010000", '1', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7639
      ("0100110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7640
      ("0000010111000111", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7641
      ("0000110111000111", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7642
      ("0000110111000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7643
      ("1000010101010100", '0', '1', "00", "101", "100", "101", '0', '-', "00"), -- i=7644
      ("1000110101010100", '1', '1', "00", "101", "100", "101", '0', '-', "00"), -- i=7645
      ("1000110101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7646
      ("1001010101010100", '0', '1', "01", "101", "100", "101", '0', '-', "00"), -- i=7647
      ("1001110101010100", '1', '1', "01", "101", "100", "101", '0', '-', "00"), -- i=7648
      ("1001110101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7649
      ("1010010101010100", '0', '1', "10", "101", "100", "101", '0', '-', "00"), -- i=7650
      ("1010110101010100", '1', '1', "10", "101", "100", "101", '0', '-', "00"), -- i=7651
      ("1010110101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7652
      ("1011010101010100", '0', '1', "11", "101", "100", "101", '0', '-', "00"), -- i=7653
      ("1011110101010100", '1', '1', "11", "101", "100", "101", '0', '-', "00"), -- i=7654
      ("1011110101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7655
      ("0101010101010000", '0', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7656
      ("0101110101010000", '1', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7657
      ("0101110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7658
      ("0100010101010000", '0', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7659
      ("0100110101010000", '1', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7660
      ("0100110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7661
      ("0000010110100000", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7662
      ("0000110110100000", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7663
      ("0000110110100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7664
      ("1000010101010101", '0', '1', "00", "101", "101", "101", '0', '-', "00"), -- i=7665
      ("1000110101010101", '1', '1', "00", "101", "101", "101", '0', '-', "00"), -- i=7666
      ("1000110101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7667
      ("1001010101010101", '0', '1', "01", "101", "101", "101", '0', '-', "00"), -- i=7668
      ("1001110101010101", '1', '1', "01", "101", "101", "101", '0', '-', "00"), -- i=7669
      ("1001110101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7670
      ("1010010101010101", '0', '1', "10", "101", "101", "101", '0', '-', "00"), -- i=7671
      ("1010110101010101", '1', '1', "10", "101", "101", "101", '0', '-', "00"), -- i=7672
      ("1010110101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7673
      ("1011010101010101", '0', '1', "11", "101", "101", "101", '0', '-', "00"), -- i=7674
      ("1011110101010101", '1', '1', "11", "101", "101", "101", '0', '-', "00"), -- i=7675
      ("1011110101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7676
      ("0101010101010000", '0', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7677
      ("0101110101010000", '1', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7678
      ("0101110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7679
      ("0100010101010000", '0', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7680
      ("0100110101010000", '1', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7681
      ("0100110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7682
      ("0000010110011011", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7683
      ("0000110110011011", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7684
      ("0000110110011011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7685
      ("1000010101010110", '0', '1', "00", "101", "110", "101", '0', '-', "00"), -- i=7686
      ("1000110101010110", '1', '1', "00", "101", "110", "101", '0', '-', "00"), -- i=7687
      ("1000110101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7688
      ("1001010101010110", '0', '1', "01", "101", "110", "101", '0', '-', "00"), -- i=7689
      ("1001110101010110", '1', '1', "01", "101", "110", "101", '0', '-', "00"), -- i=7690
      ("1001110101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7691
      ("1010010101010110", '0', '1', "10", "101", "110", "101", '0', '-', "00"), -- i=7692
      ("1010110101010110", '1', '1', "10", "101", "110", "101", '0', '-', "00"), -- i=7693
      ("1010110101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7694
      ("1011010101010110", '0', '1', "11", "101", "110", "101", '0', '-', "00"), -- i=7695
      ("1011110101010110", '1', '1', "11", "101", "110", "101", '0', '-', "00"), -- i=7696
      ("1011110101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7697
      ("0101010101010000", '0', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7698
      ("0101110101010000", '1', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7699
      ("0101110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7700
      ("0100010101010000", '0', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7701
      ("0100110101010000", '1', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7702
      ("0100110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7703
      ("0000010111001010", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7704
      ("0000110111001010", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7705
      ("0000110111001010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7706
      ("1000010101010111", '0', '1', "00", "101", "111", "101", '0', '-', "00"), -- i=7707
      ("1000110101010111", '1', '1', "00", "101", "111", "101", '0', '-', "00"), -- i=7708
      ("1000110101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7709
      ("1001010101010111", '0', '1', "01", "101", "111", "101", '0', '-', "00"), -- i=7710
      ("1001110101010111", '1', '1', "01", "101", "111", "101", '0', '-', "00"), -- i=7711
      ("1001110101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7712
      ("1010010101010111", '0', '1', "10", "101", "111", "101", '0', '-', "00"), -- i=7713
      ("1010110101010111", '1', '1', "10", "101", "111", "101", '0', '-', "00"), -- i=7714
      ("1010110101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7715
      ("1011010101010111", '0', '1', "11", "101", "111", "101", '0', '-', "00"), -- i=7716
      ("1011110101010111", '1', '1', "11", "101", "111", "101", '0', '-', "00"), -- i=7717
      ("1011110101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7718
      ("0101010101010000", '0', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7719
      ("0101110101010000", '1', '1', "--", "101", "---", "101", '0', '1', "01"), -- i=7720
      ("0101110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7721
      ("0100010101010000", '0', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7722
      ("0100110101010000", '1', '0', "--", "101", "101", "---", '1', '-', "--"), -- i=7723
      ("0100110101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7724
      ("0000010111011000", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7725
      ("0000110111011000", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7726
      ("0000110111011000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7727
      ("1000010101100000", '0', '1', "00", "110", "000", "101", '0', '-', "00"), -- i=7728
      ("1000110101100000", '1', '1', "00", "110", "000", "101", '0', '-', "00"), -- i=7729
      ("1000110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7730
      ("1001010101100000", '0', '1', "01", "110", "000", "101", '0', '-', "00"), -- i=7731
      ("1001110101100000", '1', '1', "01", "110", "000", "101", '0', '-', "00"), -- i=7732
      ("1001110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7733
      ("1010010101100000", '0', '1', "10", "110", "000", "101", '0', '-', "00"), -- i=7734
      ("1010110101100000", '1', '1', "10", "110", "000", "101", '0', '-', "00"), -- i=7735
      ("1010110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7736
      ("1011010101100000", '0', '1', "11", "110", "000", "101", '0', '-', "00"), -- i=7737
      ("1011110101100000", '1', '1', "11", "110", "000", "101", '0', '-', "00"), -- i=7738
      ("1011110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7739
      ("0101010101100000", '0', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7740
      ("0101110101100000", '1', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7741
      ("0101110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7742
      ("0100010101100000", '0', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7743
      ("0100110101100000", '1', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7744
      ("0100110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7745
      ("0000010110110010", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7746
      ("0000110110110010", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7747
      ("0000110110110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7748
      ("1000010101100001", '0', '1', "00", "110", "001", "101", '0', '-', "00"), -- i=7749
      ("1000110101100001", '1', '1', "00", "110", "001", "101", '0', '-', "00"), -- i=7750
      ("1000110101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7751
      ("1001010101100001", '0', '1', "01", "110", "001", "101", '0', '-', "00"), -- i=7752
      ("1001110101100001", '1', '1', "01", "110", "001", "101", '0', '-', "00"), -- i=7753
      ("1001110101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7754
      ("1010010101100001", '0', '1', "10", "110", "001", "101", '0', '-', "00"), -- i=7755
      ("1010110101100001", '1', '1', "10", "110", "001", "101", '0', '-', "00"), -- i=7756
      ("1010110101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7757
      ("1011010101100001", '0', '1', "11", "110", "001", "101", '0', '-', "00"), -- i=7758
      ("1011110101100001", '1', '1', "11", "110", "001", "101", '0', '-', "00"), -- i=7759
      ("1011110101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7760
      ("0101010101100000", '0', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7761
      ("0101110101100000", '1', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7762
      ("0101110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7763
      ("0100010101100000", '0', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7764
      ("0100110101100000", '1', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7765
      ("0100110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7766
      ("0000010100011011", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7767
      ("0000110100011011", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7768
      ("0000110100011011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7769
      ("1000010101100010", '0', '1', "00", "110", "010", "101", '0', '-', "00"), -- i=7770
      ("1000110101100010", '1', '1', "00", "110", "010", "101", '0', '-', "00"), -- i=7771
      ("1000110101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7772
      ("1001010101100010", '0', '1', "01", "110", "010", "101", '0', '-', "00"), -- i=7773
      ("1001110101100010", '1', '1', "01", "110", "010", "101", '0', '-', "00"), -- i=7774
      ("1001110101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7775
      ("1010010101100010", '0', '1', "10", "110", "010", "101", '0', '-', "00"), -- i=7776
      ("1010110101100010", '1', '1', "10", "110", "010", "101", '0', '-', "00"), -- i=7777
      ("1010110101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7778
      ("1011010101100010", '0', '1', "11", "110", "010", "101", '0', '-', "00"), -- i=7779
      ("1011110101100010", '1', '1', "11", "110", "010", "101", '0', '-', "00"), -- i=7780
      ("1011110101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7781
      ("0101010101100000", '0', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7782
      ("0101110101100000", '1', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7783
      ("0101110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7784
      ("0100010101100000", '0', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7785
      ("0100110101100000", '1', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7786
      ("0100110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7787
      ("0000010100010000", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7788
      ("0000110100010000", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7789
      ("0000110100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7790
      ("1000010101100011", '0', '1', "00", "110", "011", "101", '0', '-', "00"), -- i=7791
      ("1000110101100011", '1', '1', "00", "110", "011", "101", '0', '-', "00"), -- i=7792
      ("1000110101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7793
      ("1001010101100011", '0', '1', "01", "110", "011", "101", '0', '-', "00"), -- i=7794
      ("1001110101100011", '1', '1', "01", "110", "011", "101", '0', '-', "00"), -- i=7795
      ("1001110101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7796
      ("1010010101100011", '0', '1', "10", "110", "011", "101", '0', '-', "00"), -- i=7797
      ("1010110101100011", '1', '1', "10", "110", "011", "101", '0', '-', "00"), -- i=7798
      ("1010110101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7799
      ("1011010101100011", '0', '1', "11", "110", "011", "101", '0', '-', "00"), -- i=7800
      ("1011110101100011", '1', '1', "11", "110", "011", "101", '0', '-', "00"), -- i=7801
      ("1011110101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7802
      ("0101010101100000", '0', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7803
      ("0101110101100000", '1', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7804
      ("0101110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7805
      ("0100010101100000", '0', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7806
      ("0100110101100000", '1', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7807
      ("0100110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7808
      ("0000010100110111", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7809
      ("0000110100110111", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7810
      ("0000110100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7811
      ("1000010101100100", '0', '1', "00", "110", "100", "101", '0', '-', "00"), -- i=7812
      ("1000110101100100", '1', '1', "00", "110", "100", "101", '0', '-', "00"), -- i=7813
      ("1000110101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7814
      ("1001010101100100", '0', '1', "01", "110", "100", "101", '0', '-', "00"), -- i=7815
      ("1001110101100100", '1', '1', "01", "110", "100", "101", '0', '-', "00"), -- i=7816
      ("1001110101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7817
      ("1010010101100100", '0', '1', "10", "110", "100", "101", '0', '-', "00"), -- i=7818
      ("1010110101100100", '1', '1', "10", "110", "100", "101", '0', '-', "00"), -- i=7819
      ("1010110101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7820
      ("1011010101100100", '0', '1', "11", "110", "100", "101", '0', '-', "00"), -- i=7821
      ("1011110101100100", '1', '1', "11", "110", "100", "101", '0', '-', "00"), -- i=7822
      ("1011110101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7823
      ("0101010101100000", '0', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7824
      ("0101110101100000", '1', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7825
      ("0101110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7826
      ("0100010101100000", '0', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7827
      ("0100110101100000", '1', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7828
      ("0100110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7829
      ("0000010110001101", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7830
      ("0000110110001101", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7831
      ("0000110110001101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7832
      ("1000010101100101", '0', '1', "00", "110", "101", "101", '0', '-', "00"), -- i=7833
      ("1000110101100101", '1', '1', "00", "110", "101", "101", '0', '-', "00"), -- i=7834
      ("1000110101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7835
      ("1001010101100101", '0', '1', "01", "110", "101", "101", '0', '-', "00"), -- i=7836
      ("1001110101100101", '1', '1', "01", "110", "101", "101", '0', '-', "00"), -- i=7837
      ("1001110101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7838
      ("1010010101100101", '0', '1', "10", "110", "101", "101", '0', '-', "00"), -- i=7839
      ("1010110101100101", '1', '1', "10", "110", "101", "101", '0', '-', "00"), -- i=7840
      ("1010110101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7841
      ("1011010101100101", '0', '1', "11", "110", "101", "101", '0', '-', "00"), -- i=7842
      ("1011110101100101", '1', '1', "11", "110", "101", "101", '0', '-', "00"), -- i=7843
      ("1011110101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7844
      ("0101010101100000", '0', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7845
      ("0101110101100000", '1', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7846
      ("0101110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7847
      ("0100010101100000", '0', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7848
      ("0100110101100000", '1', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7849
      ("0100110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7850
      ("0000010111010110", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7851
      ("0000110111010110", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7852
      ("0000110111010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7853
      ("1000010101100110", '0', '1', "00", "110", "110", "101", '0', '-', "00"), -- i=7854
      ("1000110101100110", '1', '1', "00", "110", "110", "101", '0', '-', "00"), -- i=7855
      ("1000110101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7856
      ("1001010101100110", '0', '1', "01", "110", "110", "101", '0', '-', "00"), -- i=7857
      ("1001110101100110", '1', '1', "01", "110", "110", "101", '0', '-', "00"), -- i=7858
      ("1001110101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7859
      ("1010010101100110", '0', '1', "10", "110", "110", "101", '0', '-', "00"), -- i=7860
      ("1010110101100110", '1', '1', "10", "110", "110", "101", '0', '-', "00"), -- i=7861
      ("1010110101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7862
      ("1011010101100110", '0', '1', "11", "110", "110", "101", '0', '-', "00"), -- i=7863
      ("1011110101100110", '1', '1', "11", "110", "110", "101", '0', '-', "00"), -- i=7864
      ("1011110101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7865
      ("0101010101100000", '0', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7866
      ("0101110101100000", '1', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7867
      ("0101110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7868
      ("0100010101100000", '0', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7869
      ("0100110101100000", '1', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7870
      ("0100110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7871
      ("0000010100011111", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7872
      ("0000110100011111", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7873
      ("0000110100011111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7874
      ("1000010101100111", '0', '1', "00", "110", "111", "101", '0', '-', "00"), -- i=7875
      ("1000110101100111", '1', '1', "00", "110", "111", "101", '0', '-', "00"), -- i=7876
      ("1000110101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7877
      ("1001010101100111", '0', '1', "01", "110", "111", "101", '0', '-', "00"), -- i=7878
      ("1001110101100111", '1', '1', "01", "110", "111", "101", '0', '-', "00"), -- i=7879
      ("1001110101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7880
      ("1010010101100111", '0', '1', "10", "110", "111", "101", '0', '-', "00"), -- i=7881
      ("1010110101100111", '1', '1', "10", "110", "111", "101", '0', '-', "00"), -- i=7882
      ("1010110101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7883
      ("1011010101100111", '0', '1', "11", "110", "111", "101", '0', '-', "00"), -- i=7884
      ("1011110101100111", '1', '1', "11", "110", "111", "101", '0', '-', "00"), -- i=7885
      ("1011110101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7886
      ("0101010101100000", '0', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7887
      ("0101110101100000", '1', '1', "--", "110", "---", "101", '0', '1', "01"), -- i=7888
      ("0101110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7889
      ("0100010101100000", '0', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7890
      ("0100110101100000", '1', '0', "--", "110", "101", "---", '1', '-', "--"), -- i=7891
      ("0100110101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7892
      ("0000010100001101", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7893
      ("0000110100001101", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7894
      ("0000110100001101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7895
      ("1000010101110000", '0', '1', "00", "111", "000", "101", '0', '-', "00"), -- i=7896
      ("1000110101110000", '1', '1', "00", "111", "000", "101", '0', '-', "00"), -- i=7897
      ("1000110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7898
      ("1001010101110000", '0', '1', "01", "111", "000", "101", '0', '-', "00"), -- i=7899
      ("1001110101110000", '1', '1', "01", "111", "000", "101", '0', '-', "00"), -- i=7900
      ("1001110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7901
      ("1010010101110000", '0', '1', "10", "111", "000", "101", '0', '-', "00"), -- i=7902
      ("1010110101110000", '1', '1', "10", "111", "000", "101", '0', '-', "00"), -- i=7903
      ("1010110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7904
      ("1011010101110000", '0', '1', "11", "111", "000", "101", '0', '-', "00"), -- i=7905
      ("1011110101110000", '1', '1', "11", "111", "000", "101", '0', '-', "00"), -- i=7906
      ("1011110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7907
      ("0101010101110000", '0', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=7908
      ("0101110101110000", '1', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=7909
      ("0101110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7910
      ("0100010101110000", '0', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=7911
      ("0100110101110000", '1', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=7912
      ("0100110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7913
      ("0000010110110001", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7914
      ("0000110110110001", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7915
      ("0000110110110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7916
      ("1000010101110001", '0', '1', "00", "111", "001", "101", '0', '-', "00"), -- i=7917
      ("1000110101110001", '1', '1', "00", "111", "001", "101", '0', '-', "00"), -- i=7918
      ("1000110101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7919
      ("1001010101110001", '0', '1', "01", "111", "001", "101", '0', '-', "00"), -- i=7920
      ("1001110101110001", '1', '1', "01", "111", "001", "101", '0', '-', "00"), -- i=7921
      ("1001110101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7922
      ("1010010101110001", '0', '1', "10", "111", "001", "101", '0', '-', "00"), -- i=7923
      ("1010110101110001", '1', '1', "10", "111", "001", "101", '0', '-', "00"), -- i=7924
      ("1010110101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7925
      ("1011010101110001", '0', '1', "11", "111", "001", "101", '0', '-', "00"), -- i=7926
      ("1011110101110001", '1', '1', "11", "111", "001", "101", '0', '-', "00"), -- i=7927
      ("1011110101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7928
      ("0101010101110000", '0', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=7929
      ("0101110101110000", '1', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=7930
      ("0101110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7931
      ("0100010101110000", '0', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=7932
      ("0100110101110000", '1', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=7933
      ("0100110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7934
      ("0000010111111110", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7935
      ("0000110111111110", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7936
      ("0000110111111110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7937
      ("1000010101110010", '0', '1', "00", "111", "010", "101", '0', '-', "00"), -- i=7938
      ("1000110101110010", '1', '1', "00", "111", "010", "101", '0', '-', "00"), -- i=7939
      ("1000110101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7940
      ("1001010101110010", '0', '1', "01", "111", "010", "101", '0', '-', "00"), -- i=7941
      ("1001110101110010", '1', '1', "01", "111", "010", "101", '0', '-', "00"), -- i=7942
      ("1001110101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7943
      ("1010010101110010", '0', '1', "10", "111", "010", "101", '0', '-', "00"), -- i=7944
      ("1010110101110010", '1', '1', "10", "111", "010", "101", '0', '-', "00"), -- i=7945
      ("1010110101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7946
      ("1011010101110010", '0', '1', "11", "111", "010", "101", '0', '-', "00"), -- i=7947
      ("1011110101110010", '1', '1', "11", "111", "010", "101", '0', '-', "00"), -- i=7948
      ("1011110101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7949
      ("0101010101110000", '0', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=7950
      ("0101110101110000", '1', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=7951
      ("0101110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7952
      ("0100010101110000", '0', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=7953
      ("0100110101110000", '1', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=7954
      ("0100110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7955
      ("0000010101000110", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7956
      ("0000110101000110", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7957
      ("0000110101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7958
      ("1000010101110011", '0', '1', "00", "111", "011", "101", '0', '-', "00"), -- i=7959
      ("1000110101110011", '1', '1', "00", "111", "011", "101", '0', '-', "00"), -- i=7960
      ("1000110101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7961
      ("1001010101110011", '0', '1', "01", "111", "011", "101", '0', '-', "00"), -- i=7962
      ("1001110101110011", '1', '1', "01", "111", "011", "101", '0', '-', "00"), -- i=7963
      ("1001110101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7964
      ("1010010101110011", '0', '1', "10", "111", "011", "101", '0', '-', "00"), -- i=7965
      ("1010110101110011", '1', '1', "10", "111", "011", "101", '0', '-', "00"), -- i=7966
      ("1010110101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7967
      ("1011010101110011", '0', '1', "11", "111", "011", "101", '0', '-', "00"), -- i=7968
      ("1011110101110011", '1', '1', "11", "111", "011", "101", '0', '-', "00"), -- i=7969
      ("1011110101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7970
      ("0101010101110000", '0', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=7971
      ("0101110101110000", '1', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=7972
      ("0101110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7973
      ("0100010101110000", '0', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=7974
      ("0100110101110000", '1', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=7975
      ("0100110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7976
      ("0000010111100010", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7977
      ("0000110111100010", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7978
      ("0000110111100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7979
      ("1000010101110100", '0', '1', "00", "111", "100", "101", '0', '-', "00"), -- i=7980
      ("1000110101110100", '1', '1', "00", "111", "100", "101", '0', '-', "00"), -- i=7981
      ("1000110101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7982
      ("1001010101110100", '0', '1', "01", "111", "100", "101", '0', '-', "00"), -- i=7983
      ("1001110101110100", '1', '1', "01", "111", "100", "101", '0', '-', "00"), -- i=7984
      ("1001110101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7985
      ("1010010101110100", '0', '1', "10", "111", "100", "101", '0', '-', "00"), -- i=7986
      ("1010110101110100", '1', '1', "10", "111", "100", "101", '0', '-', "00"), -- i=7987
      ("1010110101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7988
      ("1011010101110100", '0', '1', "11", "111", "100", "101", '0', '-', "00"), -- i=7989
      ("1011110101110100", '1', '1', "11", "111", "100", "101", '0', '-', "00"), -- i=7990
      ("1011110101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7991
      ("0101010101110000", '0', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=7992
      ("0101110101110000", '1', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=7993
      ("0101110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7994
      ("0100010101110000", '0', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=7995
      ("0100110101110000", '1', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=7996
      ("0100110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=7997
      ("0000010101111100", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7998
      ("0000110101111100", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=7999
      ("0000110101111100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8000
      ("1000010101110101", '0', '1', "00", "111", "101", "101", '0', '-', "00"), -- i=8001
      ("1000110101110101", '1', '1', "00", "111", "101", "101", '0', '-', "00"), -- i=8002
      ("1000110101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8003
      ("1001010101110101", '0', '1', "01", "111", "101", "101", '0', '-', "00"), -- i=8004
      ("1001110101110101", '1', '1', "01", "111", "101", "101", '0', '-', "00"), -- i=8005
      ("1001110101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8006
      ("1010010101110101", '0', '1', "10", "111", "101", "101", '0', '-', "00"), -- i=8007
      ("1010110101110101", '1', '1', "10", "111", "101", "101", '0', '-', "00"), -- i=8008
      ("1010110101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8009
      ("1011010101110101", '0', '1', "11", "111", "101", "101", '0', '-', "00"), -- i=8010
      ("1011110101110101", '1', '1', "11", "111", "101", "101", '0', '-', "00"), -- i=8011
      ("1011110101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8012
      ("0101010101110000", '0', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=8013
      ("0101110101110000", '1', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=8014
      ("0101110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8015
      ("0100010101110000", '0', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=8016
      ("0100110101110000", '1', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=8017
      ("0100110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8018
      ("0000010111010010", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=8019
      ("0000110111010010", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=8020
      ("0000110111010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8021
      ("1000010101110110", '0', '1', "00", "111", "110", "101", '0', '-', "00"), -- i=8022
      ("1000110101110110", '1', '1', "00", "111", "110", "101", '0', '-', "00"), -- i=8023
      ("1000110101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8024
      ("1001010101110110", '0', '1', "01", "111", "110", "101", '0', '-', "00"), -- i=8025
      ("1001110101110110", '1', '1', "01", "111", "110", "101", '0', '-', "00"), -- i=8026
      ("1001110101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8027
      ("1010010101110110", '0', '1', "10", "111", "110", "101", '0', '-', "00"), -- i=8028
      ("1010110101110110", '1', '1', "10", "111", "110", "101", '0', '-', "00"), -- i=8029
      ("1010110101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8030
      ("1011010101110110", '0', '1', "11", "111", "110", "101", '0', '-', "00"), -- i=8031
      ("1011110101110110", '1', '1', "11", "111", "110", "101", '0', '-', "00"), -- i=8032
      ("1011110101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8033
      ("0101010101110000", '0', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=8034
      ("0101110101110000", '1', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=8035
      ("0101110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8036
      ("0100010101110000", '0', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=8037
      ("0100110101110000", '1', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=8038
      ("0100110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8039
      ("0000010111010001", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=8040
      ("0000110111010001", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=8041
      ("0000110111010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8042
      ("1000010101110111", '0', '1', "00", "111", "111", "101", '0', '-', "00"), -- i=8043
      ("1000110101110111", '1', '1', "00", "111", "111", "101", '0', '-', "00"), -- i=8044
      ("1000110101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8045
      ("1001010101110111", '0', '1', "01", "111", "111", "101", '0', '-', "00"), -- i=8046
      ("1001110101110111", '1', '1', "01", "111", "111", "101", '0', '-', "00"), -- i=8047
      ("1001110101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8048
      ("1010010101110111", '0', '1', "10", "111", "111", "101", '0', '-', "00"), -- i=8049
      ("1010110101110111", '1', '1', "10", "111", "111", "101", '0', '-', "00"), -- i=8050
      ("1010110101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8051
      ("1011010101110111", '0', '1', "11", "111", "111", "101", '0', '-', "00"), -- i=8052
      ("1011110101110111", '1', '1', "11", "111", "111", "101", '0', '-', "00"), -- i=8053
      ("1011110101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8054
      ("0101010101110000", '0', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=8055
      ("0101110101110000", '1', '1', "--", "111", "---", "101", '0', '1', "01"), -- i=8056
      ("0101110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8057
      ("0100010101110000", '0', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=8058
      ("0100110101110000", '1', '0', "--", "111", "101", "---", '1', '-', "--"), -- i=8059
      ("0100110101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8060
      ("0000010100000010", '0', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=8061
      ("0000110100000010", '1', '1', "--", "---", "---", "101", '0', '-', "10"), -- i=8062
      ("0000110100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8063
      ("1000011000000000", '0', '1', "00", "000", "000", "110", '0', '-', "00"), -- i=8064
      ("1000111000000000", '1', '1', "00", "000", "000", "110", '0', '-', "00"), -- i=8065
      ("1000111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8066
      ("1001011000000000", '0', '1', "01", "000", "000", "110", '0', '-', "00"), -- i=8067
      ("1001111000000000", '1', '1', "01", "000", "000", "110", '0', '-', "00"), -- i=8068
      ("1001111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8069
      ("1010011000000000", '0', '1', "10", "000", "000", "110", '0', '-', "00"), -- i=8070
      ("1010111000000000", '1', '1', "10", "000", "000", "110", '0', '-', "00"), -- i=8071
      ("1010111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8072
      ("1011011000000000", '0', '1', "11", "000", "000", "110", '0', '-', "00"), -- i=8073
      ("1011111000000000", '1', '1', "11", "000", "000", "110", '0', '-', "00"), -- i=8074
      ("1011111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8075
      ("0101011000000000", '0', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8076
      ("0101111000000000", '1', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8077
      ("0101111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8078
      ("0100011000000000", '0', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8079
      ("0100111000000000", '1', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8080
      ("0100111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8081
      ("0000011011011011", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8082
      ("0000111011011011", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8083
      ("0000111011011011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8084
      ("1000011000000001", '0', '1', "00", "000", "001", "110", '0', '-', "00"), -- i=8085
      ("1000111000000001", '1', '1', "00", "000", "001", "110", '0', '-', "00"), -- i=8086
      ("1000111000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8087
      ("1001011000000001", '0', '1', "01", "000", "001", "110", '0', '-', "00"), -- i=8088
      ("1001111000000001", '1', '1', "01", "000", "001", "110", '0', '-', "00"), -- i=8089
      ("1001111000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8090
      ("1010011000000001", '0', '1', "10", "000", "001", "110", '0', '-', "00"), -- i=8091
      ("1010111000000001", '1', '1', "10", "000", "001", "110", '0', '-', "00"), -- i=8092
      ("1010111000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8093
      ("1011011000000001", '0', '1', "11", "000", "001", "110", '0', '-', "00"), -- i=8094
      ("1011111000000001", '1', '1', "11", "000", "001", "110", '0', '-', "00"), -- i=8095
      ("1011111000000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8096
      ("0101011000000000", '0', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8097
      ("0101111000000000", '1', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8098
      ("0101111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8099
      ("0100011000000000", '0', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8100
      ("0100111000000000", '1', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8101
      ("0100111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8102
      ("0000011010110110", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8103
      ("0000111010110110", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8104
      ("0000111010110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8105
      ("1000011000000010", '0', '1', "00", "000", "010", "110", '0', '-', "00"), -- i=8106
      ("1000111000000010", '1', '1', "00", "000", "010", "110", '0', '-', "00"), -- i=8107
      ("1000111000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8108
      ("1001011000000010", '0', '1', "01", "000", "010", "110", '0', '-', "00"), -- i=8109
      ("1001111000000010", '1', '1', "01", "000", "010", "110", '0', '-', "00"), -- i=8110
      ("1001111000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8111
      ("1010011000000010", '0', '1', "10", "000", "010", "110", '0', '-', "00"), -- i=8112
      ("1010111000000010", '1', '1', "10", "000", "010", "110", '0', '-', "00"), -- i=8113
      ("1010111000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8114
      ("1011011000000010", '0', '1', "11", "000", "010", "110", '0', '-', "00"), -- i=8115
      ("1011111000000010", '1', '1', "11", "000", "010", "110", '0', '-', "00"), -- i=8116
      ("1011111000000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8117
      ("0101011000000000", '0', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8118
      ("0101111000000000", '1', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8119
      ("0101111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8120
      ("0100011000000000", '0', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8121
      ("0100111000000000", '1', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8122
      ("0100111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8123
      ("0000011011100110", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8124
      ("0000111011100110", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8125
      ("0000111011100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8126
      ("1000011000000011", '0', '1', "00", "000", "011", "110", '0', '-', "00"), -- i=8127
      ("1000111000000011", '1', '1', "00", "000", "011", "110", '0', '-', "00"), -- i=8128
      ("1000111000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8129
      ("1001011000000011", '0', '1', "01", "000", "011", "110", '0', '-', "00"), -- i=8130
      ("1001111000000011", '1', '1', "01", "000", "011", "110", '0', '-', "00"), -- i=8131
      ("1001111000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8132
      ("1010011000000011", '0', '1', "10", "000", "011", "110", '0', '-', "00"), -- i=8133
      ("1010111000000011", '1', '1', "10", "000", "011", "110", '0', '-', "00"), -- i=8134
      ("1010111000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8135
      ("1011011000000011", '0', '1', "11", "000", "011", "110", '0', '-', "00"), -- i=8136
      ("1011111000000011", '1', '1', "11", "000", "011", "110", '0', '-', "00"), -- i=8137
      ("1011111000000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8138
      ("0101011000000000", '0', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8139
      ("0101111000000000", '1', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8140
      ("0101111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8141
      ("0100011000000000", '0', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8142
      ("0100111000000000", '1', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8143
      ("0100111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8144
      ("0000011010001000", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8145
      ("0000111010001000", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8146
      ("0000111010001000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8147
      ("1000011000000100", '0', '1', "00", "000", "100", "110", '0', '-', "00"), -- i=8148
      ("1000111000000100", '1', '1', "00", "000", "100", "110", '0', '-', "00"), -- i=8149
      ("1000111000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8150
      ("1001011000000100", '0', '1', "01", "000", "100", "110", '0', '-', "00"), -- i=8151
      ("1001111000000100", '1', '1', "01", "000", "100", "110", '0', '-', "00"), -- i=8152
      ("1001111000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8153
      ("1010011000000100", '0', '1', "10", "000", "100", "110", '0', '-', "00"), -- i=8154
      ("1010111000000100", '1', '1', "10", "000", "100", "110", '0', '-', "00"), -- i=8155
      ("1010111000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8156
      ("1011011000000100", '0', '1', "11", "000", "100", "110", '0', '-', "00"), -- i=8157
      ("1011111000000100", '1', '1', "11", "000", "100", "110", '0', '-', "00"), -- i=8158
      ("1011111000000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8159
      ("0101011000000000", '0', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8160
      ("0101111000000000", '1', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8161
      ("0101111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8162
      ("0100011000000000", '0', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8163
      ("0100111000000000", '1', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8164
      ("0100111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8165
      ("0000011001000100", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8166
      ("0000111001000100", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8167
      ("0000111001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8168
      ("1000011000000101", '0', '1', "00", "000", "101", "110", '0', '-', "00"), -- i=8169
      ("1000111000000101", '1', '1', "00", "000", "101", "110", '0', '-', "00"), -- i=8170
      ("1000111000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8171
      ("1001011000000101", '0', '1', "01", "000", "101", "110", '0', '-', "00"), -- i=8172
      ("1001111000000101", '1', '1', "01", "000", "101", "110", '0', '-', "00"), -- i=8173
      ("1001111000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8174
      ("1010011000000101", '0', '1', "10", "000", "101", "110", '0', '-', "00"), -- i=8175
      ("1010111000000101", '1', '1', "10", "000", "101", "110", '0', '-', "00"), -- i=8176
      ("1010111000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8177
      ("1011011000000101", '0', '1', "11", "000", "101", "110", '0', '-', "00"), -- i=8178
      ("1011111000000101", '1', '1', "11", "000", "101", "110", '0', '-', "00"), -- i=8179
      ("1011111000000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8180
      ("0101011000000000", '0', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8181
      ("0101111000000000", '1', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8182
      ("0101111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8183
      ("0100011000000000", '0', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8184
      ("0100111000000000", '1', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8185
      ("0100111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8186
      ("0000011001101100", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8187
      ("0000111001101100", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8188
      ("0000111001101100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8189
      ("1000011000000110", '0', '1', "00", "000", "110", "110", '0', '-', "00"), -- i=8190
      ("1000111000000110", '1', '1', "00", "000", "110", "110", '0', '-', "00"), -- i=8191
      ("1000111000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8192
      ("1001011000000110", '0', '1', "01", "000", "110", "110", '0', '-', "00"), -- i=8193
      ("1001111000000110", '1', '1', "01", "000", "110", "110", '0', '-', "00"), -- i=8194
      ("1001111000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8195
      ("1010011000000110", '0', '1', "10", "000", "110", "110", '0', '-', "00"), -- i=8196
      ("1010111000000110", '1', '1', "10", "000", "110", "110", '0', '-', "00"), -- i=8197
      ("1010111000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8198
      ("1011011000000110", '0', '1', "11", "000", "110", "110", '0', '-', "00"), -- i=8199
      ("1011111000000110", '1', '1', "11", "000", "110", "110", '0', '-', "00"), -- i=8200
      ("1011111000000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8201
      ("0101011000000000", '0', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8202
      ("0101111000000000", '1', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8203
      ("0101111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8204
      ("0100011000000000", '0', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8205
      ("0100111000000000", '1', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8206
      ("0100111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8207
      ("0000011011011111", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8208
      ("0000111011011111", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8209
      ("0000111011011111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8210
      ("1000011000000111", '0', '1', "00", "000", "111", "110", '0', '-', "00"), -- i=8211
      ("1000111000000111", '1', '1', "00", "000", "111", "110", '0', '-', "00"), -- i=8212
      ("1000111000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8213
      ("1001011000000111", '0', '1', "01", "000", "111", "110", '0', '-', "00"), -- i=8214
      ("1001111000000111", '1', '1', "01", "000", "111", "110", '0', '-', "00"), -- i=8215
      ("1001111000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8216
      ("1010011000000111", '0', '1', "10", "000", "111", "110", '0', '-', "00"), -- i=8217
      ("1010111000000111", '1', '1', "10", "000", "111", "110", '0', '-', "00"), -- i=8218
      ("1010111000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8219
      ("1011011000000111", '0', '1', "11", "000", "111", "110", '0', '-', "00"), -- i=8220
      ("1011111000000111", '1', '1', "11", "000", "111", "110", '0', '-', "00"), -- i=8221
      ("1011111000000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8222
      ("0101011000000000", '0', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8223
      ("0101111000000000", '1', '1', "--", "000", "---", "110", '0', '1', "01"), -- i=8224
      ("0101111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8225
      ("0100011000000000", '0', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8226
      ("0100111000000000", '1', '0', "--", "000", "110", "---", '1', '-', "--"), -- i=8227
      ("0100111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8228
      ("0000011001000001", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8229
      ("0000111001000001", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8230
      ("0000111001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8231
      ("1000011000010000", '0', '1', "00", "001", "000", "110", '0', '-', "00"), -- i=8232
      ("1000111000010000", '1', '1', "00", "001", "000", "110", '0', '-', "00"), -- i=8233
      ("1000111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8234
      ("1001011000010000", '0', '1', "01", "001", "000", "110", '0', '-', "00"), -- i=8235
      ("1001111000010000", '1', '1', "01", "001", "000", "110", '0', '-', "00"), -- i=8236
      ("1001111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8237
      ("1010011000010000", '0', '1', "10", "001", "000", "110", '0', '-', "00"), -- i=8238
      ("1010111000010000", '1', '1', "10", "001", "000", "110", '0', '-', "00"), -- i=8239
      ("1010111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8240
      ("1011011000010000", '0', '1', "11", "001", "000", "110", '0', '-', "00"), -- i=8241
      ("1011111000010000", '1', '1', "11", "001", "000", "110", '0', '-', "00"), -- i=8242
      ("1011111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8243
      ("0101011000010000", '0', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8244
      ("0101111000010000", '1', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8245
      ("0101111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8246
      ("0100011000010000", '0', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8247
      ("0100111000010000", '1', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8248
      ("0100111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8249
      ("0000011011110001", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8250
      ("0000111011110001", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8251
      ("0000111011110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8252
      ("1000011000010001", '0', '1', "00", "001", "001", "110", '0', '-', "00"), -- i=8253
      ("1000111000010001", '1', '1', "00", "001", "001", "110", '0', '-', "00"), -- i=8254
      ("1000111000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8255
      ("1001011000010001", '0', '1', "01", "001", "001", "110", '0', '-', "00"), -- i=8256
      ("1001111000010001", '1', '1', "01", "001", "001", "110", '0', '-', "00"), -- i=8257
      ("1001111000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8258
      ("1010011000010001", '0', '1', "10", "001", "001", "110", '0', '-', "00"), -- i=8259
      ("1010111000010001", '1', '1', "10", "001", "001", "110", '0', '-', "00"), -- i=8260
      ("1010111000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8261
      ("1011011000010001", '0', '1', "11", "001", "001", "110", '0', '-', "00"), -- i=8262
      ("1011111000010001", '1', '1', "11", "001", "001", "110", '0', '-', "00"), -- i=8263
      ("1011111000010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8264
      ("0101011000010000", '0', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8265
      ("0101111000010000", '1', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8266
      ("0101111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8267
      ("0100011000010000", '0', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8268
      ("0100111000010000", '1', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8269
      ("0100111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8270
      ("0000011001001111", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8271
      ("0000111001001111", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8272
      ("0000111001001111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8273
      ("1000011000010010", '0', '1', "00", "001", "010", "110", '0', '-', "00"), -- i=8274
      ("1000111000010010", '1', '1', "00", "001", "010", "110", '0', '-', "00"), -- i=8275
      ("1000111000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8276
      ("1001011000010010", '0', '1', "01", "001", "010", "110", '0', '-', "00"), -- i=8277
      ("1001111000010010", '1', '1', "01", "001", "010", "110", '0', '-', "00"), -- i=8278
      ("1001111000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8279
      ("1010011000010010", '0', '1', "10", "001", "010", "110", '0', '-', "00"), -- i=8280
      ("1010111000010010", '1', '1', "10", "001", "010", "110", '0', '-', "00"), -- i=8281
      ("1010111000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8282
      ("1011011000010010", '0', '1', "11", "001", "010", "110", '0', '-', "00"), -- i=8283
      ("1011111000010010", '1', '1', "11", "001", "010", "110", '0', '-', "00"), -- i=8284
      ("1011111000010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8285
      ("0101011000010000", '0', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8286
      ("0101111000010000", '1', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8287
      ("0101111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8288
      ("0100011000010000", '0', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8289
      ("0100111000010000", '1', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8290
      ("0100111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8291
      ("0000011000001010", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8292
      ("0000111000001010", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8293
      ("0000111000001010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8294
      ("1000011000010011", '0', '1', "00", "001", "011", "110", '0', '-', "00"), -- i=8295
      ("1000111000010011", '1', '1', "00", "001", "011", "110", '0', '-', "00"), -- i=8296
      ("1000111000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8297
      ("1001011000010011", '0', '1', "01", "001", "011", "110", '0', '-', "00"), -- i=8298
      ("1001111000010011", '1', '1', "01", "001", "011", "110", '0', '-', "00"), -- i=8299
      ("1001111000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8300
      ("1010011000010011", '0', '1', "10", "001", "011", "110", '0', '-', "00"), -- i=8301
      ("1010111000010011", '1', '1', "10", "001", "011", "110", '0', '-', "00"), -- i=8302
      ("1010111000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8303
      ("1011011000010011", '0', '1', "11", "001", "011", "110", '0', '-', "00"), -- i=8304
      ("1011111000010011", '1', '1', "11", "001", "011", "110", '0', '-', "00"), -- i=8305
      ("1011111000010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8306
      ("0101011000010000", '0', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8307
      ("0101111000010000", '1', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8308
      ("0101111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8309
      ("0100011000010000", '0', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8310
      ("0100111000010000", '1', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8311
      ("0100111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8312
      ("0000011011111000", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8313
      ("0000111011111000", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8314
      ("0000111011111000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8315
      ("1000011000010100", '0', '1', "00", "001", "100", "110", '0', '-', "00"), -- i=8316
      ("1000111000010100", '1', '1', "00", "001", "100", "110", '0', '-', "00"), -- i=8317
      ("1000111000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8318
      ("1001011000010100", '0', '1', "01", "001", "100", "110", '0', '-', "00"), -- i=8319
      ("1001111000010100", '1', '1', "01", "001", "100", "110", '0', '-', "00"), -- i=8320
      ("1001111000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8321
      ("1010011000010100", '0', '1', "10", "001", "100", "110", '0', '-', "00"), -- i=8322
      ("1010111000010100", '1', '1', "10", "001", "100", "110", '0', '-', "00"), -- i=8323
      ("1010111000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8324
      ("1011011000010100", '0', '1', "11", "001", "100", "110", '0', '-', "00"), -- i=8325
      ("1011111000010100", '1', '1', "11", "001", "100", "110", '0', '-', "00"), -- i=8326
      ("1011111000010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8327
      ("0101011000010000", '0', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8328
      ("0101111000010000", '1', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8329
      ("0101111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8330
      ("0100011000010000", '0', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8331
      ("0100111000010000", '1', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8332
      ("0100111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8333
      ("0000011000000000", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8334
      ("0000111000000000", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8335
      ("0000111000000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8336
      ("1000011000010101", '0', '1', "00", "001", "101", "110", '0', '-', "00"), -- i=8337
      ("1000111000010101", '1', '1', "00", "001", "101", "110", '0', '-', "00"), -- i=8338
      ("1000111000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8339
      ("1001011000010101", '0', '1', "01", "001", "101", "110", '0', '-', "00"), -- i=8340
      ("1001111000010101", '1', '1', "01", "001", "101", "110", '0', '-', "00"), -- i=8341
      ("1001111000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8342
      ("1010011000010101", '0', '1', "10", "001", "101", "110", '0', '-', "00"), -- i=8343
      ("1010111000010101", '1', '1', "10", "001", "101", "110", '0', '-', "00"), -- i=8344
      ("1010111000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8345
      ("1011011000010101", '0', '1', "11", "001", "101", "110", '0', '-', "00"), -- i=8346
      ("1011111000010101", '1', '1', "11", "001", "101", "110", '0', '-', "00"), -- i=8347
      ("1011111000010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8348
      ("0101011000010000", '0', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8349
      ("0101111000010000", '1', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8350
      ("0101111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8351
      ("0100011000010000", '0', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8352
      ("0100111000010000", '1', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8353
      ("0100111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8354
      ("0000011011010010", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8355
      ("0000111011010010", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8356
      ("0000111011010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8357
      ("1000011000010110", '0', '1', "00", "001", "110", "110", '0', '-', "00"), -- i=8358
      ("1000111000010110", '1', '1', "00", "001", "110", "110", '0', '-', "00"), -- i=8359
      ("1000111000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8360
      ("1001011000010110", '0', '1', "01", "001", "110", "110", '0', '-', "00"), -- i=8361
      ("1001111000010110", '1', '1', "01", "001", "110", "110", '0', '-', "00"), -- i=8362
      ("1001111000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8363
      ("1010011000010110", '0', '1', "10", "001", "110", "110", '0', '-', "00"), -- i=8364
      ("1010111000010110", '1', '1', "10", "001", "110", "110", '0', '-', "00"), -- i=8365
      ("1010111000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8366
      ("1011011000010110", '0', '1', "11", "001", "110", "110", '0', '-', "00"), -- i=8367
      ("1011111000010110", '1', '1', "11", "001", "110", "110", '0', '-', "00"), -- i=8368
      ("1011111000010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8369
      ("0101011000010000", '0', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8370
      ("0101111000010000", '1', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8371
      ("0101111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8372
      ("0100011000010000", '0', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8373
      ("0100111000010000", '1', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8374
      ("0100111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8375
      ("0000011000001001", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8376
      ("0000111000001001", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8377
      ("0000111000001001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8378
      ("1000011000010111", '0', '1', "00", "001", "111", "110", '0', '-', "00"), -- i=8379
      ("1000111000010111", '1', '1', "00", "001", "111", "110", '0', '-', "00"), -- i=8380
      ("1000111000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8381
      ("1001011000010111", '0', '1', "01", "001", "111", "110", '0', '-', "00"), -- i=8382
      ("1001111000010111", '1', '1', "01", "001", "111", "110", '0', '-', "00"), -- i=8383
      ("1001111000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8384
      ("1010011000010111", '0', '1', "10", "001", "111", "110", '0', '-', "00"), -- i=8385
      ("1010111000010111", '1', '1', "10", "001", "111", "110", '0', '-', "00"), -- i=8386
      ("1010111000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8387
      ("1011011000010111", '0', '1', "11", "001", "111", "110", '0', '-', "00"), -- i=8388
      ("1011111000010111", '1', '1', "11", "001", "111", "110", '0', '-', "00"), -- i=8389
      ("1011111000010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8390
      ("0101011000010000", '0', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8391
      ("0101111000010000", '1', '1', "--", "001", "---", "110", '0', '1', "01"), -- i=8392
      ("0101111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8393
      ("0100011000010000", '0', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8394
      ("0100111000010000", '1', '0', "--", "001", "110", "---", '1', '-', "--"), -- i=8395
      ("0100111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8396
      ("0000011000101110", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8397
      ("0000111000101110", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8398
      ("0000111000101110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8399
      ("1000011000100000", '0', '1', "00", "010", "000", "110", '0', '-', "00"), -- i=8400
      ("1000111000100000", '1', '1', "00", "010", "000", "110", '0', '-', "00"), -- i=8401
      ("1000111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8402
      ("1001011000100000", '0', '1', "01", "010", "000", "110", '0', '-', "00"), -- i=8403
      ("1001111000100000", '1', '1', "01", "010", "000", "110", '0', '-', "00"), -- i=8404
      ("1001111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8405
      ("1010011000100000", '0', '1', "10", "010", "000", "110", '0', '-', "00"), -- i=8406
      ("1010111000100000", '1', '1', "10", "010", "000", "110", '0', '-', "00"), -- i=8407
      ("1010111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8408
      ("1011011000100000", '0', '1', "11", "010", "000", "110", '0', '-', "00"), -- i=8409
      ("1011111000100000", '1', '1', "11", "010", "000", "110", '0', '-', "00"), -- i=8410
      ("1011111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8411
      ("0101011000100000", '0', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8412
      ("0101111000100000", '1', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8413
      ("0101111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8414
      ("0100011000100000", '0', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8415
      ("0100111000100000", '1', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8416
      ("0100111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8417
      ("0000011000110110", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8418
      ("0000111000110110", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8419
      ("0000111000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8420
      ("1000011000100001", '0', '1', "00", "010", "001", "110", '0', '-', "00"), -- i=8421
      ("1000111000100001", '1', '1', "00", "010", "001", "110", '0', '-', "00"), -- i=8422
      ("1000111000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8423
      ("1001011000100001", '0', '1', "01", "010", "001", "110", '0', '-', "00"), -- i=8424
      ("1001111000100001", '1', '1', "01", "010", "001", "110", '0', '-', "00"), -- i=8425
      ("1001111000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8426
      ("1010011000100001", '0', '1', "10", "010", "001", "110", '0', '-', "00"), -- i=8427
      ("1010111000100001", '1', '1', "10", "010", "001", "110", '0', '-', "00"), -- i=8428
      ("1010111000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8429
      ("1011011000100001", '0', '1', "11", "010", "001", "110", '0', '-', "00"), -- i=8430
      ("1011111000100001", '1', '1', "11", "010", "001", "110", '0', '-', "00"), -- i=8431
      ("1011111000100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8432
      ("0101011000100000", '0', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8433
      ("0101111000100000", '1', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8434
      ("0101111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8435
      ("0100011000100000", '0', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8436
      ("0100111000100000", '1', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8437
      ("0100111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8438
      ("0000011001001101", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8439
      ("0000111001001101", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8440
      ("0000111001001101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8441
      ("1000011000100010", '0', '1', "00", "010", "010", "110", '0', '-', "00"), -- i=8442
      ("1000111000100010", '1', '1', "00", "010", "010", "110", '0', '-', "00"), -- i=8443
      ("1000111000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8444
      ("1001011000100010", '0', '1', "01", "010", "010", "110", '0', '-', "00"), -- i=8445
      ("1001111000100010", '1', '1', "01", "010", "010", "110", '0', '-', "00"), -- i=8446
      ("1001111000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8447
      ("1010011000100010", '0', '1', "10", "010", "010", "110", '0', '-', "00"), -- i=8448
      ("1010111000100010", '1', '1', "10", "010", "010", "110", '0', '-', "00"), -- i=8449
      ("1010111000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8450
      ("1011011000100010", '0', '1', "11", "010", "010", "110", '0', '-', "00"), -- i=8451
      ("1011111000100010", '1', '1', "11", "010", "010", "110", '0', '-', "00"), -- i=8452
      ("1011111000100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8453
      ("0101011000100000", '0', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8454
      ("0101111000100000", '1', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8455
      ("0101111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8456
      ("0100011000100000", '0', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8457
      ("0100111000100000", '1', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8458
      ("0100111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8459
      ("0000011000111110", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8460
      ("0000111000111110", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8461
      ("0000111000111110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8462
      ("1000011000100011", '0', '1', "00", "010", "011", "110", '0', '-', "00"), -- i=8463
      ("1000111000100011", '1', '1', "00", "010", "011", "110", '0', '-', "00"), -- i=8464
      ("1000111000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8465
      ("1001011000100011", '0', '1', "01", "010", "011", "110", '0', '-', "00"), -- i=8466
      ("1001111000100011", '1', '1', "01", "010", "011", "110", '0', '-', "00"), -- i=8467
      ("1001111000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8468
      ("1010011000100011", '0', '1', "10", "010", "011", "110", '0', '-', "00"), -- i=8469
      ("1010111000100011", '1', '1', "10", "010", "011", "110", '0', '-', "00"), -- i=8470
      ("1010111000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8471
      ("1011011000100011", '0', '1', "11", "010", "011", "110", '0', '-', "00"), -- i=8472
      ("1011111000100011", '1', '1', "11", "010", "011", "110", '0', '-', "00"), -- i=8473
      ("1011111000100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8474
      ("0101011000100000", '0', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8475
      ("0101111000100000", '1', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8476
      ("0101111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8477
      ("0100011000100000", '0', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8478
      ("0100111000100000", '1', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8479
      ("0100111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8480
      ("0000011010101011", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8481
      ("0000111010101011", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8482
      ("0000111010101011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8483
      ("1000011000100100", '0', '1', "00", "010", "100", "110", '0', '-', "00"), -- i=8484
      ("1000111000100100", '1', '1', "00", "010", "100", "110", '0', '-', "00"), -- i=8485
      ("1000111000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8486
      ("1001011000100100", '0', '1', "01", "010", "100", "110", '0', '-', "00"), -- i=8487
      ("1001111000100100", '1', '1', "01", "010", "100", "110", '0', '-', "00"), -- i=8488
      ("1001111000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8489
      ("1010011000100100", '0', '1', "10", "010", "100", "110", '0', '-', "00"), -- i=8490
      ("1010111000100100", '1', '1', "10", "010", "100", "110", '0', '-', "00"), -- i=8491
      ("1010111000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8492
      ("1011011000100100", '0', '1', "11", "010", "100", "110", '0', '-', "00"), -- i=8493
      ("1011111000100100", '1', '1', "11", "010", "100", "110", '0', '-', "00"), -- i=8494
      ("1011111000100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8495
      ("0101011000100000", '0', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8496
      ("0101111000100000", '1', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8497
      ("0101111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8498
      ("0100011000100000", '0', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8499
      ("0100111000100000", '1', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8500
      ("0100111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8501
      ("0000011010011001", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8502
      ("0000111010011001", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8503
      ("0000111010011001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8504
      ("1000011000100101", '0', '1', "00", "010", "101", "110", '0', '-', "00"), -- i=8505
      ("1000111000100101", '1', '1', "00", "010", "101", "110", '0', '-', "00"), -- i=8506
      ("1000111000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8507
      ("1001011000100101", '0', '1', "01", "010", "101", "110", '0', '-', "00"), -- i=8508
      ("1001111000100101", '1', '1', "01", "010", "101", "110", '0', '-', "00"), -- i=8509
      ("1001111000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8510
      ("1010011000100101", '0', '1', "10", "010", "101", "110", '0', '-', "00"), -- i=8511
      ("1010111000100101", '1', '1', "10", "010", "101", "110", '0', '-', "00"), -- i=8512
      ("1010111000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8513
      ("1011011000100101", '0', '1', "11", "010", "101", "110", '0', '-', "00"), -- i=8514
      ("1011111000100101", '1', '1', "11", "010", "101", "110", '0', '-', "00"), -- i=8515
      ("1011111000100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8516
      ("0101011000100000", '0', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8517
      ("0101111000100000", '1', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8518
      ("0101111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8519
      ("0100011000100000", '0', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8520
      ("0100111000100000", '1', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8521
      ("0100111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8522
      ("0000011001101001", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8523
      ("0000111001101001", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8524
      ("0000111001101001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8525
      ("1000011000100110", '0', '1', "00", "010", "110", "110", '0', '-', "00"), -- i=8526
      ("1000111000100110", '1', '1', "00", "010", "110", "110", '0', '-', "00"), -- i=8527
      ("1000111000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8528
      ("1001011000100110", '0', '1', "01", "010", "110", "110", '0', '-', "00"), -- i=8529
      ("1001111000100110", '1', '1', "01", "010", "110", "110", '0', '-', "00"), -- i=8530
      ("1001111000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8531
      ("1010011000100110", '0', '1', "10", "010", "110", "110", '0', '-', "00"), -- i=8532
      ("1010111000100110", '1', '1', "10", "010", "110", "110", '0', '-', "00"), -- i=8533
      ("1010111000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8534
      ("1011011000100110", '0', '1', "11", "010", "110", "110", '0', '-', "00"), -- i=8535
      ("1011111000100110", '1', '1', "11", "010", "110", "110", '0', '-', "00"), -- i=8536
      ("1011111000100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8537
      ("0101011000100000", '0', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8538
      ("0101111000100000", '1', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8539
      ("0101111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8540
      ("0100011000100000", '0', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8541
      ("0100111000100000", '1', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8542
      ("0100111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8543
      ("0000011001101100", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8544
      ("0000111001101100", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8545
      ("0000111001101100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8546
      ("1000011000100111", '0', '1', "00", "010", "111", "110", '0', '-', "00"), -- i=8547
      ("1000111000100111", '1', '1', "00", "010", "111", "110", '0', '-', "00"), -- i=8548
      ("1000111000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8549
      ("1001011000100111", '0', '1', "01", "010", "111", "110", '0', '-', "00"), -- i=8550
      ("1001111000100111", '1', '1', "01", "010", "111", "110", '0', '-', "00"), -- i=8551
      ("1001111000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8552
      ("1010011000100111", '0', '1', "10", "010", "111", "110", '0', '-', "00"), -- i=8553
      ("1010111000100111", '1', '1', "10", "010", "111", "110", '0', '-', "00"), -- i=8554
      ("1010111000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8555
      ("1011011000100111", '0', '1', "11", "010", "111", "110", '0', '-', "00"), -- i=8556
      ("1011111000100111", '1', '1', "11", "010", "111", "110", '0', '-', "00"), -- i=8557
      ("1011111000100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8558
      ("0101011000100000", '0', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8559
      ("0101111000100000", '1', '1', "--", "010", "---", "110", '0', '1', "01"), -- i=8560
      ("0101111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8561
      ("0100011000100000", '0', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8562
      ("0100111000100000", '1', '0', "--", "010", "110", "---", '1', '-', "--"), -- i=8563
      ("0100111000100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8564
      ("0000011011010110", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8565
      ("0000111011010110", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8566
      ("0000111011010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8567
      ("1000011000110000", '0', '1', "00", "011", "000", "110", '0', '-', "00"), -- i=8568
      ("1000111000110000", '1', '1', "00", "011", "000", "110", '0', '-', "00"), -- i=8569
      ("1000111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8570
      ("1001011000110000", '0', '1', "01", "011", "000", "110", '0', '-', "00"), -- i=8571
      ("1001111000110000", '1', '1', "01", "011", "000", "110", '0', '-', "00"), -- i=8572
      ("1001111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8573
      ("1010011000110000", '0', '1', "10", "011", "000", "110", '0', '-', "00"), -- i=8574
      ("1010111000110000", '1', '1', "10", "011", "000", "110", '0', '-', "00"), -- i=8575
      ("1010111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8576
      ("1011011000110000", '0', '1', "11", "011", "000", "110", '0', '-', "00"), -- i=8577
      ("1011111000110000", '1', '1', "11", "011", "000", "110", '0', '-', "00"), -- i=8578
      ("1011111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8579
      ("0101011000110000", '0', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8580
      ("0101111000110000", '1', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8581
      ("0101111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8582
      ("0100011000110000", '0', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8583
      ("0100111000110000", '1', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8584
      ("0100111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8585
      ("0000011010010111", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8586
      ("0000111010010111", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8587
      ("0000111010010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8588
      ("1000011000110001", '0', '1', "00", "011", "001", "110", '0', '-', "00"), -- i=8589
      ("1000111000110001", '1', '1', "00", "011", "001", "110", '0', '-', "00"), -- i=8590
      ("1000111000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8591
      ("1001011000110001", '0', '1', "01", "011", "001", "110", '0', '-', "00"), -- i=8592
      ("1001111000110001", '1', '1', "01", "011", "001", "110", '0', '-', "00"), -- i=8593
      ("1001111000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8594
      ("1010011000110001", '0', '1', "10", "011", "001", "110", '0', '-', "00"), -- i=8595
      ("1010111000110001", '1', '1', "10", "011", "001", "110", '0', '-', "00"), -- i=8596
      ("1010111000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8597
      ("1011011000110001", '0', '1', "11", "011", "001", "110", '0', '-', "00"), -- i=8598
      ("1011111000110001", '1', '1', "11", "011", "001", "110", '0', '-', "00"), -- i=8599
      ("1011111000110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8600
      ("0101011000110000", '0', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8601
      ("0101111000110000", '1', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8602
      ("0101111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8603
      ("0100011000110000", '0', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8604
      ("0100111000110000", '1', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8605
      ("0100111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8606
      ("0000011001110110", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8607
      ("0000111001110110", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8608
      ("0000111001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8609
      ("1000011000110010", '0', '1', "00", "011", "010", "110", '0', '-', "00"), -- i=8610
      ("1000111000110010", '1', '1', "00", "011", "010", "110", '0', '-', "00"), -- i=8611
      ("1000111000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8612
      ("1001011000110010", '0', '1', "01", "011", "010", "110", '0', '-', "00"), -- i=8613
      ("1001111000110010", '1', '1', "01", "011", "010", "110", '0', '-', "00"), -- i=8614
      ("1001111000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8615
      ("1010011000110010", '0', '1', "10", "011", "010", "110", '0', '-', "00"), -- i=8616
      ("1010111000110010", '1', '1', "10", "011", "010", "110", '0', '-', "00"), -- i=8617
      ("1010111000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8618
      ("1011011000110010", '0', '1', "11", "011", "010", "110", '0', '-', "00"), -- i=8619
      ("1011111000110010", '1', '1', "11", "011", "010", "110", '0', '-', "00"), -- i=8620
      ("1011111000110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8621
      ("0101011000110000", '0', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8622
      ("0101111000110000", '1', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8623
      ("0101111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8624
      ("0100011000110000", '0', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8625
      ("0100111000110000", '1', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8626
      ("0100111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8627
      ("0000011001111011", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8628
      ("0000111001111011", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8629
      ("0000111001111011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8630
      ("1000011000110011", '0', '1', "00", "011", "011", "110", '0', '-', "00"), -- i=8631
      ("1000111000110011", '1', '1', "00", "011", "011", "110", '0', '-', "00"), -- i=8632
      ("1000111000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8633
      ("1001011000110011", '0', '1', "01", "011", "011", "110", '0', '-', "00"), -- i=8634
      ("1001111000110011", '1', '1', "01", "011", "011", "110", '0', '-', "00"), -- i=8635
      ("1001111000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8636
      ("1010011000110011", '0', '1', "10", "011", "011", "110", '0', '-', "00"), -- i=8637
      ("1010111000110011", '1', '1', "10", "011", "011", "110", '0', '-', "00"), -- i=8638
      ("1010111000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8639
      ("1011011000110011", '0', '1', "11", "011", "011", "110", '0', '-', "00"), -- i=8640
      ("1011111000110011", '1', '1', "11", "011", "011", "110", '0', '-', "00"), -- i=8641
      ("1011111000110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8642
      ("0101011000110000", '0', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8643
      ("0101111000110000", '1', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8644
      ("0101111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8645
      ("0100011000110000", '0', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8646
      ("0100111000110000", '1', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8647
      ("0100111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8648
      ("0000011000111111", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8649
      ("0000111000111111", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8650
      ("0000111000111111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8651
      ("1000011000110100", '0', '1', "00", "011", "100", "110", '0', '-', "00"), -- i=8652
      ("1000111000110100", '1', '1', "00", "011", "100", "110", '0', '-', "00"), -- i=8653
      ("1000111000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8654
      ("1001011000110100", '0', '1', "01", "011", "100", "110", '0', '-', "00"), -- i=8655
      ("1001111000110100", '1', '1', "01", "011", "100", "110", '0', '-', "00"), -- i=8656
      ("1001111000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8657
      ("1010011000110100", '0', '1', "10", "011", "100", "110", '0', '-', "00"), -- i=8658
      ("1010111000110100", '1', '1', "10", "011", "100", "110", '0', '-', "00"), -- i=8659
      ("1010111000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8660
      ("1011011000110100", '0', '1', "11", "011", "100", "110", '0', '-', "00"), -- i=8661
      ("1011111000110100", '1', '1', "11", "011", "100", "110", '0', '-', "00"), -- i=8662
      ("1011111000110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8663
      ("0101011000110000", '0', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8664
      ("0101111000110000", '1', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8665
      ("0101111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8666
      ("0100011000110000", '0', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8667
      ("0100111000110000", '1', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8668
      ("0100111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8669
      ("0000011001101011", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8670
      ("0000111001101011", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8671
      ("0000111001101011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8672
      ("1000011000110101", '0', '1', "00", "011", "101", "110", '0', '-', "00"), -- i=8673
      ("1000111000110101", '1', '1', "00", "011", "101", "110", '0', '-', "00"), -- i=8674
      ("1000111000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8675
      ("1001011000110101", '0', '1', "01", "011", "101", "110", '0', '-', "00"), -- i=8676
      ("1001111000110101", '1', '1', "01", "011", "101", "110", '0', '-', "00"), -- i=8677
      ("1001111000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8678
      ("1010011000110101", '0', '1', "10", "011", "101", "110", '0', '-', "00"), -- i=8679
      ("1010111000110101", '1', '1', "10", "011", "101", "110", '0', '-', "00"), -- i=8680
      ("1010111000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8681
      ("1011011000110101", '0', '1', "11", "011", "101", "110", '0', '-', "00"), -- i=8682
      ("1011111000110101", '1', '1', "11", "011", "101", "110", '0', '-', "00"), -- i=8683
      ("1011111000110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8684
      ("0101011000110000", '0', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8685
      ("0101111000110000", '1', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8686
      ("0101111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8687
      ("0100011000110000", '0', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8688
      ("0100111000110000", '1', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8689
      ("0100111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8690
      ("0000011000111100", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8691
      ("0000111000111100", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8692
      ("0000111000111100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8693
      ("1000011000110110", '0', '1', "00", "011", "110", "110", '0', '-', "00"), -- i=8694
      ("1000111000110110", '1', '1', "00", "011", "110", "110", '0', '-', "00"), -- i=8695
      ("1000111000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8696
      ("1001011000110110", '0', '1', "01", "011", "110", "110", '0', '-', "00"), -- i=8697
      ("1001111000110110", '1', '1', "01", "011", "110", "110", '0', '-', "00"), -- i=8698
      ("1001111000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8699
      ("1010011000110110", '0', '1', "10", "011", "110", "110", '0', '-', "00"), -- i=8700
      ("1010111000110110", '1', '1', "10", "011", "110", "110", '0', '-', "00"), -- i=8701
      ("1010111000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8702
      ("1011011000110110", '0', '1', "11", "011", "110", "110", '0', '-', "00"), -- i=8703
      ("1011111000110110", '1', '1', "11", "011", "110", "110", '0', '-', "00"), -- i=8704
      ("1011111000110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8705
      ("0101011000110000", '0', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8706
      ("0101111000110000", '1', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8707
      ("0101111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8708
      ("0100011000110000", '0', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8709
      ("0100111000110000", '1', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8710
      ("0100111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8711
      ("0000011010100100", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8712
      ("0000111010100100", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8713
      ("0000111010100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8714
      ("1000011000110111", '0', '1', "00", "011", "111", "110", '0', '-', "00"), -- i=8715
      ("1000111000110111", '1', '1', "00", "011", "111", "110", '0', '-', "00"), -- i=8716
      ("1000111000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8717
      ("1001011000110111", '0', '1', "01", "011", "111", "110", '0', '-', "00"), -- i=8718
      ("1001111000110111", '1', '1', "01", "011", "111", "110", '0', '-', "00"), -- i=8719
      ("1001111000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8720
      ("1010011000110111", '0', '1', "10", "011", "111", "110", '0', '-', "00"), -- i=8721
      ("1010111000110111", '1', '1', "10", "011", "111", "110", '0', '-', "00"), -- i=8722
      ("1010111000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8723
      ("1011011000110111", '0', '1', "11", "011", "111", "110", '0', '-', "00"), -- i=8724
      ("1011111000110111", '1', '1', "11", "011", "111", "110", '0', '-', "00"), -- i=8725
      ("1011111000110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8726
      ("0101011000110000", '0', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8727
      ("0101111000110000", '1', '1', "--", "011", "---", "110", '0', '1', "01"), -- i=8728
      ("0101111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8729
      ("0100011000110000", '0', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8730
      ("0100111000110000", '1', '0', "--", "011", "110", "---", '1', '-', "--"), -- i=8731
      ("0100111000110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8732
      ("0000011001010110", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8733
      ("0000111001010110", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8734
      ("0000111001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8735
      ("1000011001000000", '0', '1', "00", "100", "000", "110", '0', '-', "00"), -- i=8736
      ("1000111001000000", '1', '1', "00", "100", "000", "110", '0', '-', "00"), -- i=8737
      ("1000111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8738
      ("1001011001000000", '0', '1', "01", "100", "000", "110", '0', '-', "00"), -- i=8739
      ("1001111001000000", '1', '1', "01", "100", "000", "110", '0', '-', "00"), -- i=8740
      ("1001111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8741
      ("1010011001000000", '0', '1', "10", "100", "000", "110", '0', '-', "00"), -- i=8742
      ("1010111001000000", '1', '1', "10", "100", "000", "110", '0', '-', "00"), -- i=8743
      ("1010111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8744
      ("1011011001000000", '0', '1', "11", "100", "000", "110", '0', '-', "00"), -- i=8745
      ("1011111001000000", '1', '1', "11", "100", "000", "110", '0', '-', "00"), -- i=8746
      ("1011111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8747
      ("0101011001000000", '0', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8748
      ("0101111001000000", '1', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8749
      ("0101111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8750
      ("0100011001000000", '0', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8751
      ("0100111001000000", '1', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8752
      ("0100111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8753
      ("0000011010110000", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8754
      ("0000111010110000", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8755
      ("0000111010110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8756
      ("1000011001000001", '0', '1', "00", "100", "001", "110", '0', '-', "00"), -- i=8757
      ("1000111001000001", '1', '1', "00", "100", "001", "110", '0', '-', "00"), -- i=8758
      ("1000111001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8759
      ("1001011001000001", '0', '1', "01", "100", "001", "110", '0', '-', "00"), -- i=8760
      ("1001111001000001", '1', '1', "01", "100", "001", "110", '0', '-', "00"), -- i=8761
      ("1001111001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8762
      ("1010011001000001", '0', '1', "10", "100", "001", "110", '0', '-', "00"), -- i=8763
      ("1010111001000001", '1', '1', "10", "100", "001", "110", '0', '-', "00"), -- i=8764
      ("1010111001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8765
      ("1011011001000001", '0', '1', "11", "100", "001", "110", '0', '-', "00"), -- i=8766
      ("1011111001000001", '1', '1', "11", "100", "001", "110", '0', '-', "00"), -- i=8767
      ("1011111001000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8768
      ("0101011001000000", '0', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8769
      ("0101111001000000", '1', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8770
      ("0101111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8771
      ("0100011001000000", '0', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8772
      ("0100111001000000", '1', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8773
      ("0100111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8774
      ("0000011011101010", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8775
      ("0000111011101010", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8776
      ("0000111011101010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8777
      ("1000011001000010", '0', '1', "00", "100", "010", "110", '0', '-', "00"), -- i=8778
      ("1000111001000010", '1', '1', "00", "100", "010", "110", '0', '-', "00"), -- i=8779
      ("1000111001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8780
      ("1001011001000010", '0', '1', "01", "100", "010", "110", '0', '-', "00"), -- i=8781
      ("1001111001000010", '1', '1', "01", "100", "010", "110", '0', '-', "00"), -- i=8782
      ("1001111001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8783
      ("1010011001000010", '0', '1', "10", "100", "010", "110", '0', '-', "00"), -- i=8784
      ("1010111001000010", '1', '1', "10", "100", "010", "110", '0', '-', "00"), -- i=8785
      ("1010111001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8786
      ("1011011001000010", '0', '1', "11", "100", "010", "110", '0', '-', "00"), -- i=8787
      ("1011111001000010", '1', '1', "11", "100", "010", "110", '0', '-', "00"), -- i=8788
      ("1011111001000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8789
      ("0101011001000000", '0', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8790
      ("0101111001000000", '1', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8791
      ("0101111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8792
      ("0100011001000000", '0', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8793
      ("0100111001000000", '1', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8794
      ("0100111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8795
      ("0000011010100000", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8796
      ("0000111010100000", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8797
      ("0000111010100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8798
      ("1000011001000011", '0', '1', "00", "100", "011", "110", '0', '-', "00"), -- i=8799
      ("1000111001000011", '1', '1', "00", "100", "011", "110", '0', '-', "00"), -- i=8800
      ("1000111001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8801
      ("1001011001000011", '0', '1', "01", "100", "011", "110", '0', '-', "00"), -- i=8802
      ("1001111001000011", '1', '1', "01", "100", "011", "110", '0', '-', "00"), -- i=8803
      ("1001111001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8804
      ("1010011001000011", '0', '1', "10", "100", "011", "110", '0', '-', "00"), -- i=8805
      ("1010111001000011", '1', '1', "10", "100", "011", "110", '0', '-', "00"), -- i=8806
      ("1010111001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8807
      ("1011011001000011", '0', '1', "11", "100", "011", "110", '0', '-', "00"), -- i=8808
      ("1011111001000011", '1', '1', "11", "100", "011", "110", '0', '-', "00"), -- i=8809
      ("1011111001000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8810
      ("0101011001000000", '0', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8811
      ("0101111001000000", '1', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8812
      ("0101111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8813
      ("0100011001000000", '0', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8814
      ("0100111001000000", '1', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8815
      ("0100111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8816
      ("0000011011010010", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8817
      ("0000111011010010", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8818
      ("0000111011010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8819
      ("1000011001000100", '0', '1', "00", "100", "100", "110", '0', '-', "00"), -- i=8820
      ("1000111001000100", '1', '1', "00", "100", "100", "110", '0', '-', "00"), -- i=8821
      ("1000111001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8822
      ("1001011001000100", '0', '1', "01", "100", "100", "110", '0', '-', "00"), -- i=8823
      ("1001111001000100", '1', '1', "01", "100", "100", "110", '0', '-', "00"), -- i=8824
      ("1001111001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8825
      ("1010011001000100", '0', '1', "10", "100", "100", "110", '0', '-', "00"), -- i=8826
      ("1010111001000100", '1', '1', "10", "100", "100", "110", '0', '-', "00"), -- i=8827
      ("1010111001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8828
      ("1011011001000100", '0', '1', "11", "100", "100", "110", '0', '-', "00"), -- i=8829
      ("1011111001000100", '1', '1', "11", "100", "100", "110", '0', '-', "00"), -- i=8830
      ("1011111001000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8831
      ("0101011001000000", '0', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8832
      ("0101111001000000", '1', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8833
      ("0101111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8834
      ("0100011001000000", '0', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8835
      ("0100111001000000", '1', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8836
      ("0100111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8837
      ("0000011001111000", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8838
      ("0000111001111000", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8839
      ("0000111001111000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8840
      ("1000011001000101", '0', '1', "00", "100", "101", "110", '0', '-', "00"), -- i=8841
      ("1000111001000101", '1', '1', "00", "100", "101", "110", '0', '-', "00"), -- i=8842
      ("1000111001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8843
      ("1001011001000101", '0', '1', "01", "100", "101", "110", '0', '-', "00"), -- i=8844
      ("1001111001000101", '1', '1', "01", "100", "101", "110", '0', '-', "00"), -- i=8845
      ("1001111001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8846
      ("1010011001000101", '0', '1', "10", "100", "101", "110", '0', '-', "00"), -- i=8847
      ("1010111001000101", '1', '1', "10", "100", "101", "110", '0', '-', "00"), -- i=8848
      ("1010111001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8849
      ("1011011001000101", '0', '1', "11", "100", "101", "110", '0', '-', "00"), -- i=8850
      ("1011111001000101", '1', '1', "11", "100", "101", "110", '0', '-', "00"), -- i=8851
      ("1011111001000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8852
      ("0101011001000000", '0', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8853
      ("0101111001000000", '1', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8854
      ("0101111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8855
      ("0100011001000000", '0', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8856
      ("0100111001000000", '1', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8857
      ("0100111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8858
      ("0000011000010000", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8859
      ("0000111000010000", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8860
      ("0000111000010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8861
      ("1000011001000110", '0', '1', "00", "100", "110", "110", '0', '-', "00"), -- i=8862
      ("1000111001000110", '1', '1', "00", "100", "110", "110", '0', '-', "00"), -- i=8863
      ("1000111001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8864
      ("1001011001000110", '0', '1', "01", "100", "110", "110", '0', '-', "00"), -- i=8865
      ("1001111001000110", '1', '1', "01", "100", "110", "110", '0', '-', "00"), -- i=8866
      ("1001111001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8867
      ("1010011001000110", '0', '1', "10", "100", "110", "110", '0', '-', "00"), -- i=8868
      ("1010111001000110", '1', '1', "10", "100", "110", "110", '0', '-', "00"), -- i=8869
      ("1010111001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8870
      ("1011011001000110", '0', '1', "11", "100", "110", "110", '0', '-', "00"), -- i=8871
      ("1011111001000110", '1', '1', "11", "100", "110", "110", '0', '-', "00"), -- i=8872
      ("1011111001000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8873
      ("0101011001000000", '0', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8874
      ("0101111001000000", '1', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8875
      ("0101111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8876
      ("0100011001000000", '0', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8877
      ("0100111001000000", '1', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8878
      ("0100111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8879
      ("0000011001011000", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8880
      ("0000111001011000", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8881
      ("0000111001011000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8882
      ("1000011001000111", '0', '1', "00", "100", "111", "110", '0', '-', "00"), -- i=8883
      ("1000111001000111", '1', '1', "00", "100", "111", "110", '0', '-', "00"), -- i=8884
      ("1000111001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8885
      ("1001011001000111", '0', '1', "01", "100", "111", "110", '0', '-', "00"), -- i=8886
      ("1001111001000111", '1', '1', "01", "100", "111", "110", '0', '-', "00"), -- i=8887
      ("1001111001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8888
      ("1010011001000111", '0', '1', "10", "100", "111", "110", '0', '-', "00"), -- i=8889
      ("1010111001000111", '1', '1', "10", "100", "111", "110", '0', '-', "00"), -- i=8890
      ("1010111001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8891
      ("1011011001000111", '0', '1', "11", "100", "111", "110", '0', '-', "00"), -- i=8892
      ("1011111001000111", '1', '1', "11", "100", "111", "110", '0', '-', "00"), -- i=8893
      ("1011111001000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8894
      ("0101011001000000", '0', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8895
      ("0101111001000000", '1', '1', "--", "100", "---", "110", '0', '1', "01"), -- i=8896
      ("0101111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8897
      ("0100011001000000", '0', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8898
      ("0100111001000000", '1', '0', "--", "100", "110", "---", '1', '-', "--"), -- i=8899
      ("0100111001000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8900
      ("0000011011111001", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8901
      ("0000111011111001", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8902
      ("0000111011111001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8903
      ("1000011001010000", '0', '1', "00", "101", "000", "110", '0', '-', "00"), -- i=8904
      ("1000111001010000", '1', '1', "00", "101", "000", "110", '0', '-', "00"), -- i=8905
      ("1000111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8906
      ("1001011001010000", '0', '1', "01", "101", "000", "110", '0', '-', "00"), -- i=8907
      ("1001111001010000", '1', '1', "01", "101", "000", "110", '0', '-', "00"), -- i=8908
      ("1001111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8909
      ("1010011001010000", '0', '1', "10", "101", "000", "110", '0', '-', "00"), -- i=8910
      ("1010111001010000", '1', '1', "10", "101", "000", "110", '0', '-', "00"), -- i=8911
      ("1010111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8912
      ("1011011001010000", '0', '1', "11", "101", "000", "110", '0', '-', "00"), -- i=8913
      ("1011111001010000", '1', '1', "11", "101", "000", "110", '0', '-', "00"), -- i=8914
      ("1011111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8915
      ("0101011001010000", '0', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=8916
      ("0101111001010000", '1', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=8917
      ("0101111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8918
      ("0100011001010000", '0', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=8919
      ("0100111001010000", '1', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=8920
      ("0100111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8921
      ("0000011000011010", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8922
      ("0000111000011010", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8923
      ("0000111000011010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8924
      ("1000011001010001", '0', '1', "00", "101", "001", "110", '0', '-', "00"), -- i=8925
      ("1000111001010001", '1', '1', "00", "101", "001", "110", '0', '-', "00"), -- i=8926
      ("1000111001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8927
      ("1001011001010001", '0', '1', "01", "101", "001", "110", '0', '-', "00"), -- i=8928
      ("1001111001010001", '1', '1', "01", "101", "001", "110", '0', '-', "00"), -- i=8929
      ("1001111001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8930
      ("1010011001010001", '0', '1', "10", "101", "001", "110", '0', '-', "00"), -- i=8931
      ("1010111001010001", '1', '1', "10", "101", "001", "110", '0', '-', "00"), -- i=8932
      ("1010111001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8933
      ("1011011001010001", '0', '1', "11", "101", "001", "110", '0', '-', "00"), -- i=8934
      ("1011111001010001", '1', '1', "11", "101", "001", "110", '0', '-', "00"), -- i=8935
      ("1011111001010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8936
      ("0101011001010000", '0', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=8937
      ("0101111001010000", '1', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=8938
      ("0101111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8939
      ("0100011001010000", '0', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=8940
      ("0100111001010000", '1', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=8941
      ("0100111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8942
      ("0000011011000000", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8943
      ("0000111011000000", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8944
      ("0000111011000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8945
      ("1000011001010010", '0', '1', "00", "101", "010", "110", '0', '-', "00"), -- i=8946
      ("1000111001010010", '1', '1', "00", "101", "010", "110", '0', '-', "00"), -- i=8947
      ("1000111001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8948
      ("1001011001010010", '0', '1', "01", "101", "010", "110", '0', '-', "00"), -- i=8949
      ("1001111001010010", '1', '1', "01", "101", "010", "110", '0', '-', "00"), -- i=8950
      ("1001111001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8951
      ("1010011001010010", '0', '1', "10", "101", "010", "110", '0', '-', "00"), -- i=8952
      ("1010111001010010", '1', '1', "10", "101", "010", "110", '0', '-', "00"), -- i=8953
      ("1010111001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8954
      ("1011011001010010", '0', '1', "11", "101", "010", "110", '0', '-', "00"), -- i=8955
      ("1011111001010010", '1', '1', "11", "101", "010", "110", '0', '-', "00"), -- i=8956
      ("1011111001010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8957
      ("0101011001010000", '0', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=8958
      ("0101111001010000", '1', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=8959
      ("0101111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8960
      ("0100011001010000", '0', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=8961
      ("0100111001010000", '1', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=8962
      ("0100111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8963
      ("0000011001101010", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8964
      ("0000111001101010", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8965
      ("0000111001101010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8966
      ("1000011001010011", '0', '1', "00", "101", "011", "110", '0', '-', "00"), -- i=8967
      ("1000111001010011", '1', '1', "00", "101", "011", "110", '0', '-', "00"), -- i=8968
      ("1000111001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8969
      ("1001011001010011", '0', '1', "01", "101", "011", "110", '0', '-', "00"), -- i=8970
      ("1001111001010011", '1', '1', "01", "101", "011", "110", '0', '-', "00"), -- i=8971
      ("1001111001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8972
      ("1010011001010011", '0', '1', "10", "101", "011", "110", '0', '-', "00"), -- i=8973
      ("1010111001010011", '1', '1', "10", "101", "011", "110", '0', '-', "00"), -- i=8974
      ("1010111001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8975
      ("1011011001010011", '0', '1', "11", "101", "011", "110", '0', '-', "00"), -- i=8976
      ("1011111001010011", '1', '1', "11", "101", "011", "110", '0', '-', "00"), -- i=8977
      ("1011111001010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8978
      ("0101011001010000", '0', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=8979
      ("0101111001010000", '1', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=8980
      ("0101111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8981
      ("0100011001010000", '0', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=8982
      ("0100111001010000", '1', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=8983
      ("0100111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8984
      ("0000011001111111", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8985
      ("0000111001111111", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=8986
      ("0000111001111111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8987
      ("1000011001010100", '0', '1', "00", "101", "100", "110", '0', '-', "00"), -- i=8988
      ("1000111001010100", '1', '1', "00", "101", "100", "110", '0', '-', "00"), -- i=8989
      ("1000111001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8990
      ("1001011001010100", '0', '1', "01", "101", "100", "110", '0', '-', "00"), -- i=8991
      ("1001111001010100", '1', '1', "01", "101", "100", "110", '0', '-', "00"), -- i=8992
      ("1001111001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8993
      ("1010011001010100", '0', '1', "10", "101", "100", "110", '0', '-', "00"), -- i=8994
      ("1010111001010100", '1', '1', "10", "101", "100", "110", '0', '-', "00"), -- i=8995
      ("1010111001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8996
      ("1011011001010100", '0', '1', "11", "101", "100", "110", '0', '-', "00"), -- i=8997
      ("1011111001010100", '1', '1', "11", "101", "100", "110", '0', '-', "00"), -- i=8998
      ("1011111001010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=8999
      ("0101011001010000", '0', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=9000
      ("0101111001010000", '1', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=9001
      ("0101111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9002
      ("0100011001010000", '0', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=9003
      ("0100111001010000", '1', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=9004
      ("0100111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9005
      ("0000011011010111", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9006
      ("0000111011010111", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9007
      ("0000111011010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9008
      ("1000011001010101", '0', '1', "00", "101", "101", "110", '0', '-', "00"), -- i=9009
      ("1000111001010101", '1', '1', "00", "101", "101", "110", '0', '-', "00"), -- i=9010
      ("1000111001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9011
      ("1001011001010101", '0', '1', "01", "101", "101", "110", '0', '-', "00"), -- i=9012
      ("1001111001010101", '1', '1', "01", "101", "101", "110", '0', '-', "00"), -- i=9013
      ("1001111001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9014
      ("1010011001010101", '0', '1', "10", "101", "101", "110", '0', '-', "00"), -- i=9015
      ("1010111001010101", '1', '1', "10", "101", "101", "110", '0', '-', "00"), -- i=9016
      ("1010111001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9017
      ("1011011001010101", '0', '1', "11", "101", "101", "110", '0', '-', "00"), -- i=9018
      ("1011111001010101", '1', '1', "11", "101", "101", "110", '0', '-', "00"), -- i=9019
      ("1011111001010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9020
      ("0101011001010000", '0', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=9021
      ("0101111001010000", '1', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=9022
      ("0101111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9023
      ("0100011001010000", '0', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=9024
      ("0100111001010000", '1', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=9025
      ("0100111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9026
      ("0000011001011001", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9027
      ("0000111001011001", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9028
      ("0000111001011001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9029
      ("1000011001010110", '0', '1', "00", "101", "110", "110", '0', '-', "00"), -- i=9030
      ("1000111001010110", '1', '1', "00", "101", "110", "110", '0', '-', "00"), -- i=9031
      ("1000111001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9032
      ("1001011001010110", '0', '1', "01", "101", "110", "110", '0', '-', "00"), -- i=9033
      ("1001111001010110", '1', '1', "01", "101", "110", "110", '0', '-', "00"), -- i=9034
      ("1001111001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9035
      ("1010011001010110", '0', '1', "10", "101", "110", "110", '0', '-', "00"), -- i=9036
      ("1010111001010110", '1', '1', "10", "101", "110", "110", '0', '-', "00"), -- i=9037
      ("1010111001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9038
      ("1011011001010110", '0', '1', "11", "101", "110", "110", '0', '-', "00"), -- i=9039
      ("1011111001010110", '1', '1', "11", "101", "110", "110", '0', '-', "00"), -- i=9040
      ("1011111001010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9041
      ("0101011001010000", '0', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=9042
      ("0101111001010000", '1', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=9043
      ("0101111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9044
      ("0100011001010000", '0', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=9045
      ("0100111001010000", '1', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=9046
      ("0100111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9047
      ("0000011001110011", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9048
      ("0000111001110011", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9049
      ("0000111001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9050
      ("1000011001010111", '0', '1', "00", "101", "111", "110", '0', '-', "00"), -- i=9051
      ("1000111001010111", '1', '1', "00", "101", "111", "110", '0', '-', "00"), -- i=9052
      ("1000111001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9053
      ("1001011001010111", '0', '1', "01", "101", "111", "110", '0', '-', "00"), -- i=9054
      ("1001111001010111", '1', '1', "01", "101", "111", "110", '0', '-', "00"), -- i=9055
      ("1001111001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9056
      ("1010011001010111", '0', '1', "10", "101", "111", "110", '0', '-', "00"), -- i=9057
      ("1010111001010111", '1', '1', "10", "101", "111", "110", '0', '-', "00"), -- i=9058
      ("1010111001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9059
      ("1011011001010111", '0', '1', "11", "101", "111", "110", '0', '-', "00"), -- i=9060
      ("1011111001010111", '1', '1', "11", "101", "111", "110", '0', '-', "00"), -- i=9061
      ("1011111001010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9062
      ("0101011001010000", '0', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=9063
      ("0101111001010000", '1', '1', "--", "101", "---", "110", '0', '1', "01"), -- i=9064
      ("0101111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9065
      ("0100011001010000", '0', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=9066
      ("0100111001010000", '1', '0', "--", "101", "110", "---", '1', '-', "--"), -- i=9067
      ("0100111001010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9068
      ("0000011001111010", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9069
      ("0000111001111010", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9070
      ("0000111001111010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9071
      ("1000011001100000", '0', '1', "00", "110", "000", "110", '0', '-', "00"), -- i=9072
      ("1000111001100000", '1', '1', "00", "110", "000", "110", '0', '-', "00"), -- i=9073
      ("1000111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9074
      ("1001011001100000", '0', '1', "01", "110", "000", "110", '0', '-', "00"), -- i=9075
      ("1001111001100000", '1', '1', "01", "110", "000", "110", '0', '-', "00"), -- i=9076
      ("1001111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9077
      ("1010011001100000", '0', '1', "10", "110", "000", "110", '0', '-', "00"), -- i=9078
      ("1010111001100000", '1', '1', "10", "110", "000", "110", '0', '-', "00"), -- i=9079
      ("1010111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9080
      ("1011011001100000", '0', '1', "11", "110", "000", "110", '0', '-', "00"), -- i=9081
      ("1011111001100000", '1', '1', "11", "110", "000", "110", '0', '-', "00"), -- i=9082
      ("1011111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9083
      ("0101011001100000", '0', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9084
      ("0101111001100000", '1', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9085
      ("0101111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9086
      ("0100011001100000", '0', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9087
      ("0100111001100000", '1', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9088
      ("0100111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9089
      ("0000011011101111", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9090
      ("0000111011101111", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9091
      ("0000111011101111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9092
      ("1000011001100001", '0', '1', "00", "110", "001", "110", '0', '-', "00"), -- i=9093
      ("1000111001100001", '1', '1', "00", "110", "001", "110", '0', '-', "00"), -- i=9094
      ("1000111001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9095
      ("1001011001100001", '0', '1', "01", "110", "001", "110", '0', '-', "00"), -- i=9096
      ("1001111001100001", '1', '1', "01", "110", "001", "110", '0', '-', "00"), -- i=9097
      ("1001111001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9098
      ("1010011001100001", '0', '1', "10", "110", "001", "110", '0', '-', "00"), -- i=9099
      ("1010111001100001", '1', '1', "10", "110", "001", "110", '0', '-', "00"), -- i=9100
      ("1010111001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9101
      ("1011011001100001", '0', '1', "11", "110", "001", "110", '0', '-', "00"), -- i=9102
      ("1011111001100001", '1', '1', "11", "110", "001", "110", '0', '-', "00"), -- i=9103
      ("1011111001100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9104
      ("0101011001100000", '0', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9105
      ("0101111001100000", '1', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9106
      ("0101111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9107
      ("0100011001100000", '0', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9108
      ("0100111001100000", '1', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9109
      ("0100111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9110
      ("0000011010000100", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9111
      ("0000111010000100", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9112
      ("0000111010000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9113
      ("1000011001100010", '0', '1', "00", "110", "010", "110", '0', '-', "00"), -- i=9114
      ("1000111001100010", '1', '1', "00", "110", "010", "110", '0', '-', "00"), -- i=9115
      ("1000111001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9116
      ("1001011001100010", '0', '1', "01", "110", "010", "110", '0', '-', "00"), -- i=9117
      ("1001111001100010", '1', '1', "01", "110", "010", "110", '0', '-', "00"), -- i=9118
      ("1001111001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9119
      ("1010011001100010", '0', '1', "10", "110", "010", "110", '0', '-', "00"), -- i=9120
      ("1010111001100010", '1', '1', "10", "110", "010", "110", '0', '-', "00"), -- i=9121
      ("1010111001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9122
      ("1011011001100010", '0', '1', "11", "110", "010", "110", '0', '-', "00"), -- i=9123
      ("1011111001100010", '1', '1', "11", "110", "010", "110", '0', '-', "00"), -- i=9124
      ("1011111001100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9125
      ("0101011001100000", '0', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9126
      ("0101111001100000", '1', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9127
      ("0101111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9128
      ("0100011001100000", '0', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9129
      ("0100111001100000", '1', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9130
      ("0100111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9131
      ("0000011001001001", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9132
      ("0000111001001001", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9133
      ("0000111001001001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9134
      ("1000011001100011", '0', '1', "00", "110", "011", "110", '0', '-', "00"), -- i=9135
      ("1000111001100011", '1', '1', "00", "110", "011", "110", '0', '-', "00"), -- i=9136
      ("1000111001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9137
      ("1001011001100011", '0', '1', "01", "110", "011", "110", '0', '-', "00"), -- i=9138
      ("1001111001100011", '1', '1', "01", "110", "011", "110", '0', '-', "00"), -- i=9139
      ("1001111001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9140
      ("1010011001100011", '0', '1', "10", "110", "011", "110", '0', '-', "00"), -- i=9141
      ("1010111001100011", '1', '1', "10", "110", "011", "110", '0', '-', "00"), -- i=9142
      ("1010111001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9143
      ("1011011001100011", '0', '1', "11", "110", "011", "110", '0', '-', "00"), -- i=9144
      ("1011111001100011", '1', '1', "11", "110", "011", "110", '0', '-', "00"), -- i=9145
      ("1011111001100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9146
      ("0101011001100000", '0', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9147
      ("0101111001100000", '1', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9148
      ("0101111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9149
      ("0100011001100000", '0', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9150
      ("0100111001100000", '1', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9151
      ("0100111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9152
      ("0000011010000101", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9153
      ("0000111010000101", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9154
      ("0000111010000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9155
      ("1000011001100100", '0', '1', "00", "110", "100", "110", '0', '-', "00"), -- i=9156
      ("1000111001100100", '1', '1', "00", "110", "100", "110", '0', '-', "00"), -- i=9157
      ("1000111001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9158
      ("1001011001100100", '0', '1', "01", "110", "100", "110", '0', '-', "00"), -- i=9159
      ("1001111001100100", '1', '1', "01", "110", "100", "110", '0', '-', "00"), -- i=9160
      ("1001111001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9161
      ("1010011001100100", '0', '1', "10", "110", "100", "110", '0', '-', "00"), -- i=9162
      ("1010111001100100", '1', '1', "10", "110", "100", "110", '0', '-', "00"), -- i=9163
      ("1010111001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9164
      ("1011011001100100", '0', '1', "11", "110", "100", "110", '0', '-', "00"), -- i=9165
      ("1011111001100100", '1', '1', "11", "110", "100", "110", '0', '-', "00"), -- i=9166
      ("1011111001100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9167
      ("0101011001100000", '0', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9168
      ("0101111001100000", '1', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9169
      ("0101111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9170
      ("0100011001100000", '0', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9171
      ("0100111001100000", '1', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9172
      ("0100111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9173
      ("0000011000111111", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9174
      ("0000111000111111", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9175
      ("0000111000111111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9176
      ("1000011001100101", '0', '1', "00", "110", "101", "110", '0', '-', "00"), -- i=9177
      ("1000111001100101", '1', '1', "00", "110", "101", "110", '0', '-', "00"), -- i=9178
      ("1000111001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9179
      ("1001011001100101", '0', '1', "01", "110", "101", "110", '0', '-', "00"), -- i=9180
      ("1001111001100101", '1', '1', "01", "110", "101", "110", '0', '-', "00"), -- i=9181
      ("1001111001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9182
      ("1010011001100101", '0', '1', "10", "110", "101", "110", '0', '-', "00"), -- i=9183
      ("1010111001100101", '1', '1', "10", "110", "101", "110", '0', '-', "00"), -- i=9184
      ("1010111001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9185
      ("1011011001100101", '0', '1', "11", "110", "101", "110", '0', '-', "00"), -- i=9186
      ("1011111001100101", '1', '1', "11", "110", "101", "110", '0', '-', "00"), -- i=9187
      ("1011111001100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9188
      ("0101011001100000", '0', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9189
      ("0101111001100000", '1', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9190
      ("0101111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9191
      ("0100011001100000", '0', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9192
      ("0100111001100000", '1', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9193
      ("0100111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9194
      ("0000011010110111", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9195
      ("0000111010110111", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9196
      ("0000111010110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9197
      ("1000011001100110", '0', '1', "00", "110", "110", "110", '0', '-', "00"), -- i=9198
      ("1000111001100110", '1', '1', "00", "110", "110", "110", '0', '-', "00"), -- i=9199
      ("1000111001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9200
      ("1001011001100110", '0', '1', "01", "110", "110", "110", '0', '-', "00"), -- i=9201
      ("1001111001100110", '1', '1', "01", "110", "110", "110", '0', '-', "00"), -- i=9202
      ("1001111001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9203
      ("1010011001100110", '0', '1', "10", "110", "110", "110", '0', '-', "00"), -- i=9204
      ("1010111001100110", '1', '1', "10", "110", "110", "110", '0', '-', "00"), -- i=9205
      ("1010111001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9206
      ("1011011001100110", '0', '1', "11", "110", "110", "110", '0', '-', "00"), -- i=9207
      ("1011111001100110", '1', '1', "11", "110", "110", "110", '0', '-', "00"), -- i=9208
      ("1011111001100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9209
      ("0101011001100000", '0', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9210
      ("0101111001100000", '1', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9211
      ("0101111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9212
      ("0100011001100000", '0', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9213
      ("0100111001100000", '1', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9214
      ("0100111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9215
      ("0000011010001001", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9216
      ("0000111010001001", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9217
      ("0000111010001001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9218
      ("1000011001100111", '0', '1', "00", "110", "111", "110", '0', '-', "00"), -- i=9219
      ("1000111001100111", '1', '1', "00", "110", "111", "110", '0', '-', "00"), -- i=9220
      ("1000111001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9221
      ("1001011001100111", '0', '1', "01", "110", "111", "110", '0', '-', "00"), -- i=9222
      ("1001111001100111", '1', '1', "01", "110", "111", "110", '0', '-', "00"), -- i=9223
      ("1001111001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9224
      ("1010011001100111", '0', '1', "10", "110", "111", "110", '0', '-', "00"), -- i=9225
      ("1010111001100111", '1', '1', "10", "110", "111", "110", '0', '-', "00"), -- i=9226
      ("1010111001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9227
      ("1011011001100111", '0', '1', "11", "110", "111", "110", '0', '-', "00"), -- i=9228
      ("1011111001100111", '1', '1', "11", "110", "111", "110", '0', '-', "00"), -- i=9229
      ("1011111001100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9230
      ("0101011001100000", '0', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9231
      ("0101111001100000", '1', '1', "--", "110", "---", "110", '0', '1', "01"), -- i=9232
      ("0101111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9233
      ("0100011001100000", '0', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9234
      ("0100111001100000", '1', '0', "--", "110", "110", "---", '1', '-', "--"), -- i=9235
      ("0100111001100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9236
      ("0000011011111000", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9237
      ("0000111011111000", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9238
      ("0000111011111000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9239
      ("1000011001110000", '0', '1', "00", "111", "000", "110", '0', '-', "00"), -- i=9240
      ("1000111001110000", '1', '1', "00", "111", "000", "110", '0', '-', "00"), -- i=9241
      ("1000111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9242
      ("1001011001110000", '0', '1', "01", "111", "000", "110", '0', '-', "00"), -- i=9243
      ("1001111001110000", '1', '1', "01", "111", "000", "110", '0', '-', "00"), -- i=9244
      ("1001111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9245
      ("1010011001110000", '0', '1', "10", "111", "000", "110", '0', '-', "00"), -- i=9246
      ("1010111001110000", '1', '1', "10", "111", "000", "110", '0', '-', "00"), -- i=9247
      ("1010111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9248
      ("1011011001110000", '0', '1', "11", "111", "000", "110", '0', '-', "00"), -- i=9249
      ("1011111001110000", '1', '1', "11", "111", "000", "110", '0', '-', "00"), -- i=9250
      ("1011111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9251
      ("0101011001110000", '0', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9252
      ("0101111001110000", '1', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9253
      ("0101111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9254
      ("0100011001110000", '0', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9255
      ("0100111001110000", '1', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9256
      ("0100111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9257
      ("0000011001101110", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9258
      ("0000111001101110", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9259
      ("0000111001101110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9260
      ("1000011001110001", '0', '1', "00", "111", "001", "110", '0', '-', "00"), -- i=9261
      ("1000111001110001", '1', '1', "00", "111", "001", "110", '0', '-', "00"), -- i=9262
      ("1000111001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9263
      ("1001011001110001", '0', '1', "01", "111", "001", "110", '0', '-', "00"), -- i=9264
      ("1001111001110001", '1', '1', "01", "111", "001", "110", '0', '-', "00"), -- i=9265
      ("1001111001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9266
      ("1010011001110001", '0', '1', "10", "111", "001", "110", '0', '-', "00"), -- i=9267
      ("1010111001110001", '1', '1', "10", "111", "001", "110", '0', '-', "00"), -- i=9268
      ("1010111001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9269
      ("1011011001110001", '0', '1', "11", "111", "001", "110", '0', '-', "00"), -- i=9270
      ("1011111001110001", '1', '1', "11", "111", "001", "110", '0', '-', "00"), -- i=9271
      ("1011111001110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9272
      ("0101011001110000", '0', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9273
      ("0101111001110000", '1', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9274
      ("0101111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9275
      ("0100011001110000", '0', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9276
      ("0100111001110000", '1', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9277
      ("0100111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9278
      ("0000011001011101", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9279
      ("0000111001011101", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9280
      ("0000111001011101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9281
      ("1000011001110010", '0', '1', "00", "111", "010", "110", '0', '-', "00"), -- i=9282
      ("1000111001110010", '1', '1', "00", "111", "010", "110", '0', '-', "00"), -- i=9283
      ("1000111001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9284
      ("1001011001110010", '0', '1', "01", "111", "010", "110", '0', '-', "00"), -- i=9285
      ("1001111001110010", '1', '1', "01", "111", "010", "110", '0', '-', "00"), -- i=9286
      ("1001111001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9287
      ("1010011001110010", '0', '1', "10", "111", "010", "110", '0', '-', "00"), -- i=9288
      ("1010111001110010", '1', '1', "10", "111", "010", "110", '0', '-', "00"), -- i=9289
      ("1010111001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9290
      ("1011011001110010", '0', '1', "11", "111", "010", "110", '0', '-', "00"), -- i=9291
      ("1011111001110010", '1', '1', "11", "111", "010", "110", '0', '-', "00"), -- i=9292
      ("1011111001110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9293
      ("0101011001110000", '0', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9294
      ("0101111001110000", '1', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9295
      ("0101111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9296
      ("0100011001110000", '0', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9297
      ("0100111001110000", '1', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9298
      ("0100111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9299
      ("0000011010111101", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9300
      ("0000111010111101", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9301
      ("0000111010111101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9302
      ("1000011001110011", '0', '1', "00", "111", "011", "110", '0', '-', "00"), -- i=9303
      ("1000111001110011", '1', '1', "00", "111", "011", "110", '0', '-', "00"), -- i=9304
      ("1000111001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9305
      ("1001011001110011", '0', '1', "01", "111", "011", "110", '0', '-', "00"), -- i=9306
      ("1001111001110011", '1', '1', "01", "111", "011", "110", '0', '-', "00"), -- i=9307
      ("1001111001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9308
      ("1010011001110011", '0', '1', "10", "111", "011", "110", '0', '-', "00"), -- i=9309
      ("1010111001110011", '1', '1', "10", "111", "011", "110", '0', '-', "00"), -- i=9310
      ("1010111001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9311
      ("1011011001110011", '0', '1', "11", "111", "011", "110", '0', '-', "00"), -- i=9312
      ("1011111001110011", '1', '1', "11", "111", "011", "110", '0', '-', "00"), -- i=9313
      ("1011111001110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9314
      ("0101011001110000", '0', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9315
      ("0101111001110000", '1', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9316
      ("0101111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9317
      ("0100011001110000", '0', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9318
      ("0100111001110000", '1', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9319
      ("0100111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9320
      ("0000011011001010", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9321
      ("0000111011001010", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9322
      ("0000111011001010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9323
      ("1000011001110100", '0', '1', "00", "111", "100", "110", '0', '-', "00"), -- i=9324
      ("1000111001110100", '1', '1', "00", "111", "100", "110", '0', '-', "00"), -- i=9325
      ("1000111001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9326
      ("1001011001110100", '0', '1', "01", "111", "100", "110", '0', '-', "00"), -- i=9327
      ("1001111001110100", '1', '1', "01", "111", "100", "110", '0', '-', "00"), -- i=9328
      ("1001111001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9329
      ("1010011001110100", '0', '1', "10", "111", "100", "110", '0', '-', "00"), -- i=9330
      ("1010111001110100", '1', '1', "10", "111", "100", "110", '0', '-', "00"), -- i=9331
      ("1010111001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9332
      ("1011011001110100", '0', '1', "11", "111", "100", "110", '0', '-', "00"), -- i=9333
      ("1011111001110100", '1', '1', "11", "111", "100", "110", '0', '-', "00"), -- i=9334
      ("1011111001110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9335
      ("0101011001110000", '0', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9336
      ("0101111001110000", '1', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9337
      ("0101111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9338
      ("0100011001110000", '0', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9339
      ("0100111001110000", '1', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9340
      ("0100111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9341
      ("0000011011100010", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9342
      ("0000111011100010", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9343
      ("0000111011100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9344
      ("1000011001110101", '0', '1', "00", "111", "101", "110", '0', '-', "00"), -- i=9345
      ("1000111001110101", '1', '1', "00", "111", "101", "110", '0', '-', "00"), -- i=9346
      ("1000111001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9347
      ("1001011001110101", '0', '1', "01", "111", "101", "110", '0', '-', "00"), -- i=9348
      ("1001111001110101", '1', '1', "01", "111", "101", "110", '0', '-', "00"), -- i=9349
      ("1001111001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9350
      ("1010011001110101", '0', '1', "10", "111", "101", "110", '0', '-', "00"), -- i=9351
      ("1010111001110101", '1', '1', "10", "111", "101", "110", '0', '-', "00"), -- i=9352
      ("1010111001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9353
      ("1011011001110101", '0', '1', "11", "111", "101", "110", '0', '-', "00"), -- i=9354
      ("1011111001110101", '1', '1', "11", "111", "101", "110", '0', '-', "00"), -- i=9355
      ("1011111001110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9356
      ("0101011001110000", '0', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9357
      ("0101111001110000", '1', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9358
      ("0101111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9359
      ("0100011001110000", '0', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9360
      ("0100111001110000", '1', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9361
      ("0100111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9362
      ("0000011010111111", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9363
      ("0000111010111111", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9364
      ("0000111010111111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9365
      ("1000011001110110", '0', '1', "00", "111", "110", "110", '0', '-', "00"), -- i=9366
      ("1000111001110110", '1', '1', "00", "111", "110", "110", '0', '-', "00"), -- i=9367
      ("1000111001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9368
      ("1001011001110110", '0', '1', "01", "111", "110", "110", '0', '-', "00"), -- i=9369
      ("1001111001110110", '1', '1', "01", "111", "110", "110", '0', '-', "00"), -- i=9370
      ("1001111001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9371
      ("1010011001110110", '0', '1', "10", "111", "110", "110", '0', '-', "00"), -- i=9372
      ("1010111001110110", '1', '1', "10", "111", "110", "110", '0', '-', "00"), -- i=9373
      ("1010111001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9374
      ("1011011001110110", '0', '1', "11", "111", "110", "110", '0', '-', "00"), -- i=9375
      ("1011111001110110", '1', '1', "11", "111", "110", "110", '0', '-', "00"), -- i=9376
      ("1011111001110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9377
      ("0101011001110000", '0', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9378
      ("0101111001110000", '1', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9379
      ("0101111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9380
      ("0100011001110000", '0', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9381
      ("0100111001110000", '1', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9382
      ("0100111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9383
      ("0000011000001110", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9384
      ("0000111000001110", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9385
      ("0000111000001110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9386
      ("1000011001110111", '0', '1', "00", "111", "111", "110", '0', '-', "00"), -- i=9387
      ("1000111001110111", '1', '1', "00", "111", "111", "110", '0', '-', "00"), -- i=9388
      ("1000111001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9389
      ("1001011001110111", '0', '1', "01", "111", "111", "110", '0', '-', "00"), -- i=9390
      ("1001111001110111", '1', '1', "01", "111", "111", "110", '0', '-', "00"), -- i=9391
      ("1001111001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9392
      ("1010011001110111", '0', '1', "10", "111", "111", "110", '0', '-', "00"), -- i=9393
      ("1010111001110111", '1', '1', "10", "111", "111", "110", '0', '-', "00"), -- i=9394
      ("1010111001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9395
      ("1011011001110111", '0', '1', "11", "111", "111", "110", '0', '-', "00"), -- i=9396
      ("1011111001110111", '1', '1', "11", "111", "111", "110", '0', '-', "00"), -- i=9397
      ("1011111001110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9398
      ("0101011001110000", '0', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9399
      ("0101111001110000", '1', '1', "--", "111", "---", "110", '0', '1', "01"), -- i=9400
      ("0101111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9401
      ("0100011001110000", '0', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9402
      ("0100111001110000", '1', '0', "--", "111", "110", "---", '1', '-', "--"), -- i=9403
      ("0100111001110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9404
      ("0000011010010000", '0', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9405
      ("0000111010010000", '1', '1', "--", "---", "---", "110", '0', '-', "10"), -- i=9406
      ("0000111010010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9407
      ("1000011100000000", '0', '1', "00", "000", "000", "111", '0', '-', "00"), -- i=9408
      ("1000111100000000", '1', '1', "00", "000", "000", "111", '0', '-', "00"), -- i=9409
      ("1000111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9410
      ("1001011100000000", '0', '1', "01", "000", "000", "111", '0', '-', "00"), -- i=9411
      ("1001111100000000", '1', '1', "01", "000", "000", "111", '0', '-', "00"), -- i=9412
      ("1001111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9413
      ("1010011100000000", '0', '1', "10", "000", "000", "111", '0', '-', "00"), -- i=9414
      ("1010111100000000", '1', '1', "10", "000", "000", "111", '0', '-', "00"), -- i=9415
      ("1010111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9416
      ("1011011100000000", '0', '1', "11", "000", "000", "111", '0', '-', "00"), -- i=9417
      ("1011111100000000", '1', '1', "11", "000", "000", "111", '0', '-', "00"), -- i=9418
      ("1011111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9419
      ("0101011100000000", '0', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9420
      ("0101111100000000", '1', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9421
      ("0101111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9422
      ("0100011100000000", '0', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9423
      ("0100111100000000", '1', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9424
      ("0100111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9425
      ("0000011100011110", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9426
      ("0000111100011110", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9427
      ("0000111100011110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9428
      ("1000011100000001", '0', '1', "00", "000", "001", "111", '0', '-', "00"), -- i=9429
      ("1000111100000001", '1', '1', "00", "000", "001", "111", '0', '-', "00"), -- i=9430
      ("1000111100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9431
      ("1001011100000001", '0', '1', "01", "000", "001", "111", '0', '-', "00"), -- i=9432
      ("1001111100000001", '1', '1', "01", "000", "001", "111", '0', '-', "00"), -- i=9433
      ("1001111100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9434
      ("1010011100000001", '0', '1', "10", "000", "001", "111", '0', '-', "00"), -- i=9435
      ("1010111100000001", '1', '1', "10", "000", "001", "111", '0', '-', "00"), -- i=9436
      ("1010111100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9437
      ("1011011100000001", '0', '1', "11", "000", "001", "111", '0', '-', "00"), -- i=9438
      ("1011111100000001", '1', '1', "11", "000", "001", "111", '0', '-', "00"), -- i=9439
      ("1011111100000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9440
      ("0101011100000000", '0', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9441
      ("0101111100000000", '1', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9442
      ("0101111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9443
      ("0100011100000000", '0', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9444
      ("0100111100000000", '1', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9445
      ("0100111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9446
      ("0000011110111100", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9447
      ("0000111110111100", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9448
      ("0000111110111100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9449
      ("1000011100000010", '0', '1', "00", "000", "010", "111", '0', '-', "00"), -- i=9450
      ("1000111100000010", '1', '1', "00", "000", "010", "111", '0', '-', "00"), -- i=9451
      ("1000111100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9452
      ("1001011100000010", '0', '1', "01", "000", "010", "111", '0', '-', "00"), -- i=9453
      ("1001111100000010", '1', '1', "01", "000", "010", "111", '0', '-', "00"), -- i=9454
      ("1001111100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9455
      ("1010011100000010", '0', '1', "10", "000", "010", "111", '0', '-', "00"), -- i=9456
      ("1010111100000010", '1', '1', "10", "000", "010", "111", '0', '-', "00"), -- i=9457
      ("1010111100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9458
      ("1011011100000010", '0', '1', "11", "000", "010", "111", '0', '-', "00"), -- i=9459
      ("1011111100000010", '1', '1', "11", "000", "010", "111", '0', '-', "00"), -- i=9460
      ("1011111100000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9461
      ("0101011100000000", '0', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9462
      ("0101111100000000", '1', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9463
      ("0101111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9464
      ("0100011100000000", '0', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9465
      ("0100111100000000", '1', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9466
      ("0100111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9467
      ("0000011111110000", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9468
      ("0000111111110000", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9469
      ("0000111111110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9470
      ("1000011100000011", '0', '1', "00", "000", "011", "111", '0', '-', "00"), -- i=9471
      ("1000111100000011", '1', '1', "00", "000", "011", "111", '0', '-', "00"), -- i=9472
      ("1000111100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9473
      ("1001011100000011", '0', '1', "01", "000", "011", "111", '0', '-', "00"), -- i=9474
      ("1001111100000011", '1', '1', "01", "000", "011", "111", '0', '-', "00"), -- i=9475
      ("1001111100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9476
      ("1010011100000011", '0', '1', "10", "000", "011", "111", '0', '-', "00"), -- i=9477
      ("1010111100000011", '1', '1', "10", "000", "011", "111", '0', '-', "00"), -- i=9478
      ("1010111100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9479
      ("1011011100000011", '0', '1', "11", "000", "011", "111", '0', '-', "00"), -- i=9480
      ("1011111100000011", '1', '1', "11", "000", "011", "111", '0', '-', "00"), -- i=9481
      ("1011111100000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9482
      ("0101011100000000", '0', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9483
      ("0101111100000000", '1', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9484
      ("0101111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9485
      ("0100011100000000", '0', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9486
      ("0100111100000000", '1', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9487
      ("0100111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9488
      ("0000011111001101", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9489
      ("0000111111001101", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9490
      ("0000111111001101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9491
      ("1000011100000100", '0', '1', "00", "000", "100", "111", '0', '-', "00"), -- i=9492
      ("1000111100000100", '1', '1', "00", "000", "100", "111", '0', '-', "00"), -- i=9493
      ("1000111100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9494
      ("1001011100000100", '0', '1', "01", "000", "100", "111", '0', '-', "00"), -- i=9495
      ("1001111100000100", '1', '1', "01", "000", "100", "111", '0', '-', "00"), -- i=9496
      ("1001111100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9497
      ("1010011100000100", '0', '1', "10", "000", "100", "111", '0', '-', "00"), -- i=9498
      ("1010111100000100", '1', '1', "10", "000", "100", "111", '0', '-', "00"), -- i=9499
      ("1010111100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9500
      ("1011011100000100", '0', '1', "11", "000", "100", "111", '0', '-', "00"), -- i=9501
      ("1011111100000100", '1', '1', "11", "000", "100", "111", '0', '-', "00"), -- i=9502
      ("1011111100000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9503
      ("0101011100000000", '0', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9504
      ("0101111100000000", '1', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9505
      ("0101111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9506
      ("0100011100000000", '0', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9507
      ("0100111100000000", '1', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9508
      ("0100111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9509
      ("0000011111110010", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9510
      ("0000111111110010", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9511
      ("0000111111110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9512
      ("1000011100000101", '0', '1', "00", "000", "101", "111", '0', '-', "00"), -- i=9513
      ("1000111100000101", '1', '1', "00", "000", "101", "111", '0', '-', "00"), -- i=9514
      ("1000111100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9515
      ("1001011100000101", '0', '1', "01", "000", "101", "111", '0', '-', "00"), -- i=9516
      ("1001111100000101", '1', '1', "01", "000", "101", "111", '0', '-', "00"), -- i=9517
      ("1001111100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9518
      ("1010011100000101", '0', '1', "10", "000", "101", "111", '0', '-', "00"), -- i=9519
      ("1010111100000101", '1', '1', "10", "000", "101", "111", '0', '-', "00"), -- i=9520
      ("1010111100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9521
      ("1011011100000101", '0', '1', "11", "000", "101", "111", '0', '-', "00"), -- i=9522
      ("1011111100000101", '1', '1', "11", "000", "101", "111", '0', '-', "00"), -- i=9523
      ("1011111100000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9524
      ("0101011100000000", '0', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9525
      ("0101111100000000", '1', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9526
      ("0101111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9527
      ("0100011100000000", '0', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9528
      ("0100111100000000", '1', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9529
      ("0100111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9530
      ("0000011100100010", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9531
      ("0000111100100010", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9532
      ("0000111100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9533
      ("1000011100000110", '0', '1', "00", "000", "110", "111", '0', '-', "00"), -- i=9534
      ("1000111100000110", '1', '1', "00", "000", "110", "111", '0', '-', "00"), -- i=9535
      ("1000111100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9536
      ("1001011100000110", '0', '1', "01", "000", "110", "111", '0', '-', "00"), -- i=9537
      ("1001111100000110", '1', '1', "01", "000", "110", "111", '0', '-', "00"), -- i=9538
      ("1001111100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9539
      ("1010011100000110", '0', '1', "10", "000", "110", "111", '0', '-', "00"), -- i=9540
      ("1010111100000110", '1', '1', "10", "000", "110", "111", '0', '-', "00"), -- i=9541
      ("1010111100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9542
      ("1011011100000110", '0', '1', "11", "000", "110", "111", '0', '-', "00"), -- i=9543
      ("1011111100000110", '1', '1', "11", "000", "110", "111", '0', '-', "00"), -- i=9544
      ("1011111100000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9545
      ("0101011100000000", '0', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9546
      ("0101111100000000", '1', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9547
      ("0101111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9548
      ("0100011100000000", '0', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9549
      ("0100111100000000", '1', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9550
      ("0100111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9551
      ("0000011101101101", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9552
      ("0000111101101101", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9553
      ("0000111101101101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9554
      ("1000011100000111", '0', '1', "00", "000", "111", "111", '0', '-', "00"), -- i=9555
      ("1000111100000111", '1', '1', "00", "000", "111", "111", '0', '-', "00"), -- i=9556
      ("1000111100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9557
      ("1001011100000111", '0', '1', "01", "000", "111", "111", '0', '-', "00"), -- i=9558
      ("1001111100000111", '1', '1', "01", "000", "111", "111", '0', '-', "00"), -- i=9559
      ("1001111100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9560
      ("1010011100000111", '0', '1', "10", "000", "111", "111", '0', '-', "00"), -- i=9561
      ("1010111100000111", '1', '1', "10", "000", "111", "111", '0', '-', "00"), -- i=9562
      ("1010111100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9563
      ("1011011100000111", '0', '1', "11", "000", "111", "111", '0', '-', "00"), -- i=9564
      ("1011111100000111", '1', '1', "11", "000", "111", "111", '0', '-', "00"), -- i=9565
      ("1011111100000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9566
      ("0101011100000000", '0', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9567
      ("0101111100000000", '1', '1', "--", "000", "---", "111", '0', '1', "01"), -- i=9568
      ("0101111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9569
      ("0100011100000000", '0', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9570
      ("0100111100000000", '1', '0', "--", "000", "111", "---", '1', '-', "--"), -- i=9571
      ("0100111100000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9572
      ("0000011110101111", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9573
      ("0000111110101111", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9574
      ("0000111110101111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9575
      ("1000011100010000", '0', '1', "00", "001", "000", "111", '0', '-', "00"), -- i=9576
      ("1000111100010000", '1', '1', "00", "001", "000", "111", '0', '-', "00"), -- i=9577
      ("1000111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9578
      ("1001011100010000", '0', '1', "01", "001", "000", "111", '0', '-', "00"), -- i=9579
      ("1001111100010000", '1', '1', "01", "001", "000", "111", '0', '-', "00"), -- i=9580
      ("1001111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9581
      ("1010011100010000", '0', '1', "10", "001", "000", "111", '0', '-', "00"), -- i=9582
      ("1010111100010000", '1', '1', "10", "001", "000", "111", '0', '-', "00"), -- i=9583
      ("1010111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9584
      ("1011011100010000", '0', '1', "11", "001", "000", "111", '0', '-', "00"), -- i=9585
      ("1011111100010000", '1', '1', "11", "001", "000", "111", '0', '-', "00"), -- i=9586
      ("1011111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9587
      ("0101011100010000", '0', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9588
      ("0101111100010000", '1', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9589
      ("0101111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9590
      ("0100011100010000", '0', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9591
      ("0100111100010000", '1', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9592
      ("0100111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9593
      ("0000011111100110", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9594
      ("0000111111100110", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9595
      ("0000111111100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9596
      ("1000011100010001", '0', '1', "00", "001", "001", "111", '0', '-', "00"), -- i=9597
      ("1000111100010001", '1', '1', "00", "001", "001", "111", '0', '-', "00"), -- i=9598
      ("1000111100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9599
      ("1001011100010001", '0', '1', "01", "001", "001", "111", '0', '-', "00"), -- i=9600
      ("1001111100010001", '1', '1', "01", "001", "001", "111", '0', '-', "00"), -- i=9601
      ("1001111100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9602
      ("1010011100010001", '0', '1', "10", "001", "001", "111", '0', '-', "00"), -- i=9603
      ("1010111100010001", '1', '1', "10", "001", "001", "111", '0', '-', "00"), -- i=9604
      ("1010111100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9605
      ("1011011100010001", '0', '1', "11", "001", "001", "111", '0', '-', "00"), -- i=9606
      ("1011111100010001", '1', '1', "11", "001", "001", "111", '0', '-', "00"), -- i=9607
      ("1011111100010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9608
      ("0101011100010000", '0', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9609
      ("0101111100010000", '1', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9610
      ("0101111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9611
      ("0100011100010000", '0', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9612
      ("0100111100010000", '1', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9613
      ("0100111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9614
      ("0000011111010101", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9615
      ("0000111111010101", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9616
      ("0000111111010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9617
      ("1000011100010010", '0', '1', "00", "001", "010", "111", '0', '-', "00"), -- i=9618
      ("1000111100010010", '1', '1', "00", "001", "010", "111", '0', '-', "00"), -- i=9619
      ("1000111100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9620
      ("1001011100010010", '0', '1', "01", "001", "010", "111", '0', '-', "00"), -- i=9621
      ("1001111100010010", '1', '1', "01", "001", "010", "111", '0', '-', "00"), -- i=9622
      ("1001111100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9623
      ("1010011100010010", '0', '1', "10", "001", "010", "111", '0', '-', "00"), -- i=9624
      ("1010111100010010", '1', '1', "10", "001", "010", "111", '0', '-', "00"), -- i=9625
      ("1010111100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9626
      ("1011011100010010", '0', '1', "11", "001", "010", "111", '0', '-', "00"), -- i=9627
      ("1011111100010010", '1', '1', "11", "001", "010", "111", '0', '-', "00"), -- i=9628
      ("1011111100010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9629
      ("0101011100010000", '0', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9630
      ("0101111100010000", '1', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9631
      ("0101111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9632
      ("0100011100010000", '0', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9633
      ("0100111100010000", '1', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9634
      ("0100111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9635
      ("0000011111010000", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9636
      ("0000111111010000", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9637
      ("0000111111010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9638
      ("1000011100010011", '0', '1', "00", "001", "011", "111", '0', '-', "00"), -- i=9639
      ("1000111100010011", '1', '1', "00", "001", "011", "111", '0', '-', "00"), -- i=9640
      ("1000111100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9641
      ("1001011100010011", '0', '1', "01", "001", "011", "111", '0', '-', "00"), -- i=9642
      ("1001111100010011", '1', '1', "01", "001", "011", "111", '0', '-', "00"), -- i=9643
      ("1001111100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9644
      ("1010011100010011", '0', '1', "10", "001", "011", "111", '0', '-', "00"), -- i=9645
      ("1010111100010011", '1', '1', "10", "001", "011", "111", '0', '-', "00"), -- i=9646
      ("1010111100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9647
      ("1011011100010011", '0', '1', "11", "001", "011", "111", '0', '-', "00"), -- i=9648
      ("1011111100010011", '1', '1', "11", "001", "011", "111", '0', '-', "00"), -- i=9649
      ("1011111100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9650
      ("0101011100010000", '0', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9651
      ("0101111100010000", '1', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9652
      ("0101111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9653
      ("0100011100010000", '0', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9654
      ("0100111100010000", '1', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9655
      ("0100111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9656
      ("0000011100110100", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9657
      ("0000111100110100", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9658
      ("0000111100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9659
      ("1000011100010100", '0', '1', "00", "001", "100", "111", '0', '-', "00"), -- i=9660
      ("1000111100010100", '1', '1', "00", "001", "100", "111", '0', '-', "00"), -- i=9661
      ("1000111100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9662
      ("1001011100010100", '0', '1', "01", "001", "100", "111", '0', '-', "00"), -- i=9663
      ("1001111100010100", '1', '1', "01", "001", "100", "111", '0', '-', "00"), -- i=9664
      ("1001111100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9665
      ("1010011100010100", '0', '1', "10", "001", "100", "111", '0', '-', "00"), -- i=9666
      ("1010111100010100", '1', '1', "10", "001", "100", "111", '0', '-', "00"), -- i=9667
      ("1010111100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9668
      ("1011011100010100", '0', '1', "11", "001", "100", "111", '0', '-', "00"), -- i=9669
      ("1011111100010100", '1', '1', "11", "001", "100", "111", '0', '-', "00"), -- i=9670
      ("1011111100010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9671
      ("0101011100010000", '0', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9672
      ("0101111100010000", '1', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9673
      ("0101111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9674
      ("0100011100010000", '0', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9675
      ("0100111100010000", '1', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9676
      ("0100111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9677
      ("0000011110001001", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9678
      ("0000111110001001", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9679
      ("0000111110001001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9680
      ("1000011100010101", '0', '1', "00", "001", "101", "111", '0', '-', "00"), -- i=9681
      ("1000111100010101", '1', '1', "00", "001", "101", "111", '0', '-', "00"), -- i=9682
      ("1000111100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9683
      ("1001011100010101", '0', '1', "01", "001", "101", "111", '0', '-', "00"), -- i=9684
      ("1001111100010101", '1', '1', "01", "001", "101", "111", '0', '-', "00"), -- i=9685
      ("1001111100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9686
      ("1010011100010101", '0', '1', "10", "001", "101", "111", '0', '-', "00"), -- i=9687
      ("1010111100010101", '1', '1', "10", "001", "101", "111", '0', '-', "00"), -- i=9688
      ("1010111100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9689
      ("1011011100010101", '0', '1', "11", "001", "101", "111", '0', '-', "00"), -- i=9690
      ("1011111100010101", '1', '1', "11", "001", "101", "111", '0', '-', "00"), -- i=9691
      ("1011111100010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9692
      ("0101011100010000", '0', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9693
      ("0101111100010000", '1', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9694
      ("0101111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9695
      ("0100011100010000", '0', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9696
      ("0100111100010000", '1', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9697
      ("0100111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9698
      ("0000011110000111", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9699
      ("0000111110000111", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9700
      ("0000111110000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9701
      ("1000011100010110", '0', '1', "00", "001", "110", "111", '0', '-', "00"), -- i=9702
      ("1000111100010110", '1', '1', "00", "001", "110", "111", '0', '-', "00"), -- i=9703
      ("1000111100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9704
      ("1001011100010110", '0', '1', "01", "001", "110", "111", '0', '-', "00"), -- i=9705
      ("1001111100010110", '1', '1', "01", "001", "110", "111", '0', '-', "00"), -- i=9706
      ("1001111100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9707
      ("1010011100010110", '0', '1', "10", "001", "110", "111", '0', '-', "00"), -- i=9708
      ("1010111100010110", '1', '1', "10", "001", "110", "111", '0', '-', "00"), -- i=9709
      ("1010111100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9710
      ("1011011100010110", '0', '1', "11", "001", "110", "111", '0', '-', "00"), -- i=9711
      ("1011111100010110", '1', '1', "11", "001", "110", "111", '0', '-', "00"), -- i=9712
      ("1011111100010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9713
      ("0101011100010000", '0', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9714
      ("0101111100010000", '1', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9715
      ("0101111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9716
      ("0100011100010000", '0', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9717
      ("0100111100010000", '1', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9718
      ("0100111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9719
      ("0000011100101100", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9720
      ("0000111100101100", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9721
      ("0000111100101100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9722
      ("1000011100010111", '0', '1', "00", "001", "111", "111", '0', '-', "00"), -- i=9723
      ("1000111100010111", '1', '1', "00", "001", "111", "111", '0', '-', "00"), -- i=9724
      ("1000111100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9725
      ("1001011100010111", '0', '1', "01", "001", "111", "111", '0', '-', "00"), -- i=9726
      ("1001111100010111", '1', '1', "01", "001", "111", "111", '0', '-', "00"), -- i=9727
      ("1001111100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9728
      ("1010011100010111", '0', '1', "10", "001", "111", "111", '0', '-', "00"), -- i=9729
      ("1010111100010111", '1', '1', "10", "001", "111", "111", '0', '-', "00"), -- i=9730
      ("1010111100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9731
      ("1011011100010111", '0', '1', "11", "001", "111", "111", '0', '-', "00"), -- i=9732
      ("1011111100010111", '1', '1', "11", "001", "111", "111", '0', '-', "00"), -- i=9733
      ("1011111100010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9734
      ("0101011100010000", '0', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9735
      ("0101111100010000", '1', '1', "--", "001", "---", "111", '0', '1', "01"), -- i=9736
      ("0101111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9737
      ("0100011100010000", '0', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9738
      ("0100111100010000", '1', '0', "--", "001", "111", "---", '1', '-', "--"), -- i=9739
      ("0100111100010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9740
      ("0000011110001001", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9741
      ("0000111110001001", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9742
      ("0000111110001001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9743
      ("1000011100100000", '0', '1', "00", "010", "000", "111", '0', '-', "00"), -- i=9744
      ("1000111100100000", '1', '1', "00", "010", "000", "111", '0', '-', "00"), -- i=9745
      ("1000111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9746
      ("1001011100100000", '0', '1', "01", "010", "000", "111", '0', '-', "00"), -- i=9747
      ("1001111100100000", '1', '1', "01", "010", "000", "111", '0', '-', "00"), -- i=9748
      ("1001111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9749
      ("1010011100100000", '0', '1', "10", "010", "000", "111", '0', '-', "00"), -- i=9750
      ("1010111100100000", '1', '1', "10", "010", "000", "111", '0', '-', "00"), -- i=9751
      ("1010111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9752
      ("1011011100100000", '0', '1', "11", "010", "000", "111", '0', '-', "00"), -- i=9753
      ("1011111100100000", '1', '1', "11", "010", "000", "111", '0', '-', "00"), -- i=9754
      ("1011111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9755
      ("0101011100100000", '0', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9756
      ("0101111100100000", '1', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9757
      ("0101111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9758
      ("0100011100100000", '0', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9759
      ("0100111100100000", '1', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9760
      ("0100111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9761
      ("0000011111111100", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9762
      ("0000111111111100", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9763
      ("0000111111111100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9764
      ("1000011100100001", '0', '1', "00", "010", "001", "111", '0', '-', "00"), -- i=9765
      ("1000111100100001", '1', '1', "00", "010", "001", "111", '0', '-', "00"), -- i=9766
      ("1000111100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9767
      ("1001011100100001", '0', '1', "01", "010", "001", "111", '0', '-', "00"), -- i=9768
      ("1001111100100001", '1', '1', "01", "010", "001", "111", '0', '-', "00"), -- i=9769
      ("1001111100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9770
      ("1010011100100001", '0', '1', "10", "010", "001", "111", '0', '-', "00"), -- i=9771
      ("1010111100100001", '1', '1', "10", "010", "001", "111", '0', '-', "00"), -- i=9772
      ("1010111100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9773
      ("1011011100100001", '0', '1', "11", "010", "001", "111", '0', '-', "00"), -- i=9774
      ("1011111100100001", '1', '1', "11", "010", "001", "111", '0', '-', "00"), -- i=9775
      ("1011111100100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9776
      ("0101011100100000", '0', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9777
      ("0101111100100000", '1', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9778
      ("0101111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9779
      ("0100011100100000", '0', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9780
      ("0100111100100000", '1', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9781
      ("0100111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9782
      ("0000011100111111", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9783
      ("0000111100111111", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9784
      ("0000111100111111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9785
      ("1000011100100010", '0', '1', "00", "010", "010", "111", '0', '-', "00"), -- i=9786
      ("1000111100100010", '1', '1', "00", "010", "010", "111", '0', '-', "00"), -- i=9787
      ("1000111100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9788
      ("1001011100100010", '0', '1', "01", "010", "010", "111", '0', '-', "00"), -- i=9789
      ("1001111100100010", '1', '1', "01", "010", "010", "111", '0', '-', "00"), -- i=9790
      ("1001111100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9791
      ("1010011100100010", '0', '1', "10", "010", "010", "111", '0', '-', "00"), -- i=9792
      ("1010111100100010", '1', '1', "10", "010", "010", "111", '0', '-', "00"), -- i=9793
      ("1010111100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9794
      ("1011011100100010", '0', '1', "11", "010", "010", "111", '0', '-', "00"), -- i=9795
      ("1011111100100010", '1', '1', "11", "010", "010", "111", '0', '-', "00"), -- i=9796
      ("1011111100100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9797
      ("0101011100100000", '0', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9798
      ("0101111100100000", '1', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9799
      ("0101111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9800
      ("0100011100100000", '0', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9801
      ("0100111100100000", '1', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9802
      ("0100111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9803
      ("0000011111100000", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9804
      ("0000111111100000", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9805
      ("0000111111100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9806
      ("1000011100100011", '0', '1', "00", "010", "011", "111", '0', '-', "00"), -- i=9807
      ("1000111100100011", '1', '1', "00", "010", "011", "111", '0', '-', "00"), -- i=9808
      ("1000111100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9809
      ("1001011100100011", '0', '1', "01", "010", "011", "111", '0', '-', "00"), -- i=9810
      ("1001111100100011", '1', '1', "01", "010", "011", "111", '0', '-', "00"), -- i=9811
      ("1001111100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9812
      ("1010011100100011", '0', '1', "10", "010", "011", "111", '0', '-', "00"), -- i=9813
      ("1010111100100011", '1', '1', "10", "010", "011", "111", '0', '-', "00"), -- i=9814
      ("1010111100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9815
      ("1011011100100011", '0', '1', "11", "010", "011", "111", '0', '-', "00"), -- i=9816
      ("1011111100100011", '1', '1', "11", "010", "011", "111", '0', '-', "00"), -- i=9817
      ("1011111100100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9818
      ("0101011100100000", '0', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9819
      ("0101111100100000", '1', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9820
      ("0101111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9821
      ("0100011100100000", '0', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9822
      ("0100111100100000", '1', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9823
      ("0100111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9824
      ("0000011110010001", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9825
      ("0000111110010001", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9826
      ("0000111110010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9827
      ("1000011100100100", '0', '1', "00", "010", "100", "111", '0', '-', "00"), -- i=9828
      ("1000111100100100", '1', '1', "00", "010", "100", "111", '0', '-', "00"), -- i=9829
      ("1000111100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9830
      ("1001011100100100", '0', '1', "01", "010", "100", "111", '0', '-', "00"), -- i=9831
      ("1001111100100100", '1', '1', "01", "010", "100", "111", '0', '-', "00"), -- i=9832
      ("1001111100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9833
      ("1010011100100100", '0', '1', "10", "010", "100", "111", '0', '-', "00"), -- i=9834
      ("1010111100100100", '1', '1', "10", "010", "100", "111", '0', '-', "00"), -- i=9835
      ("1010111100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9836
      ("1011011100100100", '0', '1', "11", "010", "100", "111", '0', '-', "00"), -- i=9837
      ("1011111100100100", '1', '1', "11", "010", "100", "111", '0', '-', "00"), -- i=9838
      ("1011111100100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9839
      ("0101011100100000", '0', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9840
      ("0101111100100000", '1', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9841
      ("0101111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9842
      ("0100011100100000", '0', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9843
      ("0100111100100000", '1', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9844
      ("0100111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9845
      ("0000011111010001", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9846
      ("0000111111010001", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9847
      ("0000111111010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9848
      ("1000011100100101", '0', '1', "00", "010", "101", "111", '0', '-', "00"), -- i=9849
      ("1000111100100101", '1', '1', "00", "010", "101", "111", '0', '-', "00"), -- i=9850
      ("1000111100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9851
      ("1001011100100101", '0', '1', "01", "010", "101", "111", '0', '-', "00"), -- i=9852
      ("1001111100100101", '1', '1', "01", "010", "101", "111", '0', '-', "00"), -- i=9853
      ("1001111100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9854
      ("1010011100100101", '0', '1', "10", "010", "101", "111", '0', '-', "00"), -- i=9855
      ("1010111100100101", '1', '1', "10", "010", "101", "111", '0', '-', "00"), -- i=9856
      ("1010111100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9857
      ("1011011100100101", '0', '1', "11", "010", "101", "111", '0', '-', "00"), -- i=9858
      ("1011111100100101", '1', '1', "11", "010", "101", "111", '0', '-', "00"), -- i=9859
      ("1011111100100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9860
      ("0101011100100000", '0', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9861
      ("0101111100100000", '1', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9862
      ("0101111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9863
      ("0100011100100000", '0', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9864
      ("0100111100100000", '1', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9865
      ("0100111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9866
      ("0000011110100110", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9867
      ("0000111110100110", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9868
      ("0000111110100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9869
      ("1000011100100110", '0', '1', "00", "010", "110", "111", '0', '-', "00"), -- i=9870
      ("1000111100100110", '1', '1', "00", "010", "110", "111", '0', '-', "00"), -- i=9871
      ("1000111100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9872
      ("1001011100100110", '0', '1', "01", "010", "110", "111", '0', '-', "00"), -- i=9873
      ("1001111100100110", '1', '1', "01", "010", "110", "111", '0', '-', "00"), -- i=9874
      ("1001111100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9875
      ("1010011100100110", '0', '1', "10", "010", "110", "111", '0', '-', "00"), -- i=9876
      ("1010111100100110", '1', '1', "10", "010", "110", "111", '0', '-', "00"), -- i=9877
      ("1010111100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9878
      ("1011011100100110", '0', '1', "11", "010", "110", "111", '0', '-', "00"), -- i=9879
      ("1011111100100110", '1', '1', "11", "010", "110", "111", '0', '-', "00"), -- i=9880
      ("1011111100100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9881
      ("0101011100100000", '0', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9882
      ("0101111100100000", '1', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9883
      ("0101111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9884
      ("0100011100100000", '0', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9885
      ("0100111100100000", '1', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9886
      ("0100111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9887
      ("0000011110010111", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9888
      ("0000111110010111", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9889
      ("0000111110010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9890
      ("1000011100100111", '0', '1', "00", "010", "111", "111", '0', '-', "00"), -- i=9891
      ("1000111100100111", '1', '1', "00", "010", "111", "111", '0', '-', "00"), -- i=9892
      ("1000111100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9893
      ("1001011100100111", '0', '1', "01", "010", "111", "111", '0', '-', "00"), -- i=9894
      ("1001111100100111", '1', '1', "01", "010", "111", "111", '0', '-', "00"), -- i=9895
      ("1001111100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9896
      ("1010011100100111", '0', '1', "10", "010", "111", "111", '0', '-', "00"), -- i=9897
      ("1010111100100111", '1', '1', "10", "010", "111", "111", '0', '-', "00"), -- i=9898
      ("1010111100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9899
      ("1011011100100111", '0', '1', "11", "010", "111", "111", '0', '-', "00"), -- i=9900
      ("1011111100100111", '1', '1', "11", "010", "111", "111", '0', '-', "00"), -- i=9901
      ("1011111100100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9902
      ("0101011100100000", '0', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9903
      ("0101111100100000", '1', '1', "--", "010", "---", "111", '0', '1', "01"), -- i=9904
      ("0101111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9905
      ("0100011100100000", '0', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9906
      ("0100111100100000", '1', '0', "--", "010", "111", "---", '1', '-', "--"), -- i=9907
      ("0100111100100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9908
      ("0000011101001100", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9909
      ("0000111101001100", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9910
      ("0000111101001100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9911
      ("1000011100110000", '0', '1', "00", "011", "000", "111", '0', '-', "00"), -- i=9912
      ("1000111100110000", '1', '1', "00", "011", "000", "111", '0', '-', "00"), -- i=9913
      ("1000111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9914
      ("1001011100110000", '0', '1', "01", "011", "000", "111", '0', '-', "00"), -- i=9915
      ("1001111100110000", '1', '1', "01", "011", "000", "111", '0', '-', "00"), -- i=9916
      ("1001111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9917
      ("1010011100110000", '0', '1', "10", "011", "000", "111", '0', '-', "00"), -- i=9918
      ("1010111100110000", '1', '1', "10", "011", "000", "111", '0', '-', "00"), -- i=9919
      ("1010111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9920
      ("1011011100110000", '0', '1', "11", "011", "000", "111", '0', '-', "00"), -- i=9921
      ("1011111100110000", '1', '1', "11", "011", "000", "111", '0', '-', "00"), -- i=9922
      ("1011111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9923
      ("0101011100110000", '0', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=9924
      ("0101111100110000", '1', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=9925
      ("0101111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9926
      ("0100011100110000", '0', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=9927
      ("0100111100110000", '1', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=9928
      ("0100111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9929
      ("0000011110010010", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9930
      ("0000111110010010", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9931
      ("0000111110010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9932
      ("1000011100110001", '0', '1', "00", "011", "001", "111", '0', '-', "00"), -- i=9933
      ("1000111100110001", '1', '1', "00", "011", "001", "111", '0', '-', "00"), -- i=9934
      ("1000111100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9935
      ("1001011100110001", '0', '1', "01", "011", "001", "111", '0', '-', "00"), -- i=9936
      ("1001111100110001", '1', '1', "01", "011", "001", "111", '0', '-', "00"), -- i=9937
      ("1001111100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9938
      ("1010011100110001", '0', '1', "10", "011", "001", "111", '0', '-', "00"), -- i=9939
      ("1010111100110001", '1', '1', "10", "011", "001", "111", '0', '-', "00"), -- i=9940
      ("1010111100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9941
      ("1011011100110001", '0', '1', "11", "011", "001", "111", '0', '-', "00"), -- i=9942
      ("1011111100110001", '1', '1', "11", "011", "001", "111", '0', '-', "00"), -- i=9943
      ("1011111100110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9944
      ("0101011100110000", '0', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=9945
      ("0101111100110000", '1', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=9946
      ("0101111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9947
      ("0100011100110000", '0', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=9948
      ("0100111100110000", '1', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=9949
      ("0100111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9950
      ("0000011101111011", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9951
      ("0000111101111011", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9952
      ("0000111101111011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9953
      ("1000011100110010", '0', '1', "00", "011", "010", "111", '0', '-', "00"), -- i=9954
      ("1000111100110010", '1', '1', "00", "011", "010", "111", '0', '-', "00"), -- i=9955
      ("1000111100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9956
      ("1001011100110010", '0', '1', "01", "011", "010", "111", '0', '-', "00"), -- i=9957
      ("1001111100110010", '1', '1', "01", "011", "010", "111", '0', '-', "00"), -- i=9958
      ("1001111100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9959
      ("1010011100110010", '0', '1', "10", "011", "010", "111", '0', '-', "00"), -- i=9960
      ("1010111100110010", '1', '1', "10", "011", "010", "111", '0', '-', "00"), -- i=9961
      ("1010111100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9962
      ("1011011100110010", '0', '1', "11", "011", "010", "111", '0', '-', "00"), -- i=9963
      ("1011111100110010", '1', '1', "11", "011", "010", "111", '0', '-', "00"), -- i=9964
      ("1011111100110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9965
      ("0101011100110000", '0', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=9966
      ("0101111100110000", '1', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=9967
      ("0101111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9968
      ("0100011100110000", '0', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=9969
      ("0100111100110000", '1', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=9970
      ("0100111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9971
      ("0000011101101000", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9972
      ("0000111101101000", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9973
      ("0000111101101000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9974
      ("1000011100110011", '0', '1', "00", "011", "011", "111", '0', '-', "00"), -- i=9975
      ("1000111100110011", '1', '1', "00", "011", "011", "111", '0', '-', "00"), -- i=9976
      ("1000111100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9977
      ("1001011100110011", '0', '1', "01", "011", "011", "111", '0', '-', "00"), -- i=9978
      ("1001111100110011", '1', '1', "01", "011", "011", "111", '0', '-', "00"), -- i=9979
      ("1001111100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9980
      ("1010011100110011", '0', '1', "10", "011", "011", "111", '0', '-', "00"), -- i=9981
      ("1010111100110011", '1', '1', "10", "011", "011", "111", '0', '-', "00"), -- i=9982
      ("1010111100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9983
      ("1011011100110011", '0', '1', "11", "011", "011", "111", '0', '-', "00"), -- i=9984
      ("1011111100110011", '1', '1', "11", "011", "011", "111", '0', '-', "00"), -- i=9985
      ("1011111100110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9986
      ("0101011100110000", '0', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=9987
      ("0101111100110000", '1', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=9988
      ("0101111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9989
      ("0100011100110000", '0', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=9990
      ("0100111100110000", '1', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=9991
      ("0100111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9992
      ("0000011111111111", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9993
      ("0000111111111111", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=9994
      ("0000111111111111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9995
      ("1000011100110100", '0', '1', "00", "011", "100", "111", '0', '-', "00"), -- i=9996
      ("1000111100110100", '1', '1', "00", "011", "100", "111", '0', '-', "00"), -- i=9997
      ("1000111100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=9998
      ("1001011100110100", '0', '1', "01", "011", "100", "111", '0', '-', "00"), -- i=9999
      ("1001111100110100", '1', '1', "01", "011", "100", "111", '0', '-', "00"), -- i=10000
      ("1001111100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10001
      ("1010011100110100", '0', '1', "10", "011", "100", "111", '0', '-', "00"), -- i=10002
      ("1010111100110100", '1', '1', "10", "011", "100", "111", '0', '-', "00"), -- i=10003
      ("1010111100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10004
      ("1011011100110100", '0', '1', "11", "011", "100", "111", '0', '-', "00"), -- i=10005
      ("1011111100110100", '1', '1', "11", "011", "100", "111", '0', '-', "00"), -- i=10006
      ("1011111100110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10007
      ("0101011100110000", '0', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=10008
      ("0101111100110000", '1', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=10009
      ("0101111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10010
      ("0100011100110000", '0', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=10011
      ("0100111100110000", '1', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=10012
      ("0100111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10013
      ("0000011110011010", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10014
      ("0000111110011010", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10015
      ("0000111110011010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10016
      ("1000011100110101", '0', '1', "00", "011", "101", "111", '0', '-', "00"), -- i=10017
      ("1000111100110101", '1', '1', "00", "011", "101", "111", '0', '-', "00"), -- i=10018
      ("1000111100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10019
      ("1001011100110101", '0', '1', "01", "011", "101", "111", '0', '-', "00"), -- i=10020
      ("1001111100110101", '1', '1', "01", "011", "101", "111", '0', '-', "00"), -- i=10021
      ("1001111100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10022
      ("1010011100110101", '0', '1', "10", "011", "101", "111", '0', '-', "00"), -- i=10023
      ("1010111100110101", '1', '1', "10", "011", "101", "111", '0', '-', "00"), -- i=10024
      ("1010111100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10025
      ("1011011100110101", '0', '1', "11", "011", "101", "111", '0', '-', "00"), -- i=10026
      ("1011111100110101", '1', '1', "11", "011", "101", "111", '0', '-', "00"), -- i=10027
      ("1011111100110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10028
      ("0101011100110000", '0', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=10029
      ("0101111100110000", '1', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=10030
      ("0101111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10031
      ("0100011100110000", '0', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=10032
      ("0100111100110000", '1', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=10033
      ("0100111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10034
      ("0000011101111001", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10035
      ("0000111101111001", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10036
      ("0000111101111001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10037
      ("1000011100110110", '0', '1', "00", "011", "110", "111", '0', '-', "00"), -- i=10038
      ("1000111100110110", '1', '1', "00", "011", "110", "111", '0', '-', "00"), -- i=10039
      ("1000111100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10040
      ("1001011100110110", '0', '1', "01", "011", "110", "111", '0', '-', "00"), -- i=10041
      ("1001111100110110", '1', '1', "01", "011", "110", "111", '0', '-', "00"), -- i=10042
      ("1001111100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10043
      ("1010011100110110", '0', '1', "10", "011", "110", "111", '0', '-', "00"), -- i=10044
      ("1010111100110110", '1', '1', "10", "011", "110", "111", '0', '-', "00"), -- i=10045
      ("1010111100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10046
      ("1011011100110110", '0', '1', "11", "011", "110", "111", '0', '-', "00"), -- i=10047
      ("1011111100110110", '1', '1', "11", "011", "110", "111", '0', '-', "00"), -- i=10048
      ("1011111100110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10049
      ("0101011100110000", '0', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=10050
      ("0101111100110000", '1', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=10051
      ("0101111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10052
      ("0100011100110000", '0', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=10053
      ("0100111100110000", '1', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=10054
      ("0100111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10055
      ("0000011110101111", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10056
      ("0000111110101111", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10057
      ("0000111110101111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10058
      ("1000011100110111", '0', '1', "00", "011", "111", "111", '0', '-', "00"), -- i=10059
      ("1000111100110111", '1', '1', "00", "011", "111", "111", '0', '-', "00"), -- i=10060
      ("1000111100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10061
      ("1001011100110111", '0', '1', "01", "011", "111", "111", '0', '-', "00"), -- i=10062
      ("1001111100110111", '1', '1', "01", "011", "111", "111", '0', '-', "00"), -- i=10063
      ("1001111100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10064
      ("1010011100110111", '0', '1', "10", "011", "111", "111", '0', '-', "00"), -- i=10065
      ("1010111100110111", '1', '1', "10", "011", "111", "111", '0', '-', "00"), -- i=10066
      ("1010111100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10067
      ("1011011100110111", '0', '1', "11", "011", "111", "111", '0', '-', "00"), -- i=10068
      ("1011111100110111", '1', '1', "11", "011", "111", "111", '0', '-', "00"), -- i=10069
      ("1011111100110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10070
      ("0101011100110000", '0', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=10071
      ("0101111100110000", '1', '1', "--", "011", "---", "111", '0', '1', "01"), -- i=10072
      ("0101111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10073
      ("0100011100110000", '0', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=10074
      ("0100111100110000", '1', '0', "--", "011", "111", "---", '1', '-', "--"), -- i=10075
      ("0100111100110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10076
      ("0000011111110100", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10077
      ("0000111111110100", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10078
      ("0000111111110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10079
      ("1000011101000000", '0', '1', "00", "100", "000", "111", '0', '-', "00"), -- i=10080
      ("1000111101000000", '1', '1', "00", "100", "000", "111", '0', '-', "00"), -- i=10081
      ("1000111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10082
      ("1001011101000000", '0', '1', "01", "100", "000", "111", '0', '-', "00"), -- i=10083
      ("1001111101000000", '1', '1', "01", "100", "000", "111", '0', '-', "00"), -- i=10084
      ("1001111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10085
      ("1010011101000000", '0', '1', "10", "100", "000", "111", '0', '-', "00"), -- i=10086
      ("1010111101000000", '1', '1', "10", "100", "000", "111", '0', '-', "00"), -- i=10087
      ("1010111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10088
      ("1011011101000000", '0', '1', "11", "100", "000", "111", '0', '-', "00"), -- i=10089
      ("1011111101000000", '1', '1', "11", "100", "000", "111", '0', '-', "00"), -- i=10090
      ("1011111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10091
      ("0101011101000000", '0', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10092
      ("0101111101000000", '1', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10093
      ("0101111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10094
      ("0100011101000000", '0', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10095
      ("0100111101000000", '1', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10096
      ("0100111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10097
      ("0000011110101111", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10098
      ("0000111110101111", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10099
      ("0000111110101111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10100
      ("1000011101000001", '0', '1', "00", "100", "001", "111", '0', '-', "00"), -- i=10101
      ("1000111101000001", '1', '1', "00", "100", "001", "111", '0', '-', "00"), -- i=10102
      ("1000111101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10103
      ("1001011101000001", '0', '1', "01", "100", "001", "111", '0', '-', "00"), -- i=10104
      ("1001111101000001", '1', '1', "01", "100", "001", "111", '0', '-', "00"), -- i=10105
      ("1001111101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10106
      ("1010011101000001", '0', '1', "10", "100", "001", "111", '0', '-', "00"), -- i=10107
      ("1010111101000001", '1', '1', "10", "100", "001", "111", '0', '-', "00"), -- i=10108
      ("1010111101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10109
      ("1011011101000001", '0', '1', "11", "100", "001", "111", '0', '-', "00"), -- i=10110
      ("1011111101000001", '1', '1', "11", "100", "001", "111", '0', '-', "00"), -- i=10111
      ("1011111101000001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10112
      ("0101011101000000", '0', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10113
      ("0101111101000000", '1', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10114
      ("0101111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10115
      ("0100011101000000", '0', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10116
      ("0100111101000000", '1', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10117
      ("0100111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10118
      ("0000011101010100", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10119
      ("0000111101010100", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10120
      ("0000111101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10121
      ("1000011101000010", '0', '1', "00", "100", "010", "111", '0', '-', "00"), -- i=10122
      ("1000111101000010", '1', '1', "00", "100", "010", "111", '0', '-', "00"), -- i=10123
      ("1000111101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10124
      ("1001011101000010", '0', '1', "01", "100", "010", "111", '0', '-', "00"), -- i=10125
      ("1001111101000010", '1', '1', "01", "100", "010", "111", '0', '-', "00"), -- i=10126
      ("1001111101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10127
      ("1010011101000010", '0', '1', "10", "100", "010", "111", '0', '-', "00"), -- i=10128
      ("1010111101000010", '1', '1', "10", "100", "010", "111", '0', '-', "00"), -- i=10129
      ("1010111101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10130
      ("1011011101000010", '0', '1', "11", "100", "010", "111", '0', '-', "00"), -- i=10131
      ("1011111101000010", '1', '1', "11", "100", "010", "111", '0', '-', "00"), -- i=10132
      ("1011111101000010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10133
      ("0101011101000000", '0', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10134
      ("0101111101000000", '1', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10135
      ("0101111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10136
      ("0100011101000000", '0', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10137
      ("0100111101000000", '1', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10138
      ("0100111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10139
      ("0000011111100100", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10140
      ("0000111111100100", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10141
      ("0000111111100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10142
      ("1000011101000011", '0', '1', "00", "100", "011", "111", '0', '-', "00"), -- i=10143
      ("1000111101000011", '1', '1', "00", "100", "011", "111", '0', '-', "00"), -- i=10144
      ("1000111101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10145
      ("1001011101000011", '0', '1', "01", "100", "011", "111", '0', '-', "00"), -- i=10146
      ("1001111101000011", '1', '1', "01", "100", "011", "111", '0', '-', "00"), -- i=10147
      ("1001111101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10148
      ("1010011101000011", '0', '1', "10", "100", "011", "111", '0', '-', "00"), -- i=10149
      ("1010111101000011", '1', '1', "10", "100", "011", "111", '0', '-', "00"), -- i=10150
      ("1010111101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10151
      ("1011011101000011", '0', '1', "11", "100", "011", "111", '0', '-', "00"), -- i=10152
      ("1011111101000011", '1', '1', "11", "100", "011", "111", '0', '-', "00"), -- i=10153
      ("1011111101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10154
      ("0101011101000000", '0', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10155
      ("0101111101000000", '1', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10156
      ("0101111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10157
      ("0100011101000000", '0', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10158
      ("0100111101000000", '1', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10159
      ("0100111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10160
      ("0000011110110111", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10161
      ("0000111110110111", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10162
      ("0000111110110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10163
      ("1000011101000100", '0', '1', "00", "100", "100", "111", '0', '-', "00"), -- i=10164
      ("1000111101000100", '1', '1', "00", "100", "100", "111", '0', '-', "00"), -- i=10165
      ("1000111101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10166
      ("1001011101000100", '0', '1', "01", "100", "100", "111", '0', '-', "00"), -- i=10167
      ("1001111101000100", '1', '1', "01", "100", "100", "111", '0', '-', "00"), -- i=10168
      ("1001111101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10169
      ("1010011101000100", '0', '1', "10", "100", "100", "111", '0', '-', "00"), -- i=10170
      ("1010111101000100", '1', '1', "10", "100", "100", "111", '0', '-', "00"), -- i=10171
      ("1010111101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10172
      ("1011011101000100", '0', '1', "11", "100", "100", "111", '0', '-', "00"), -- i=10173
      ("1011111101000100", '1', '1', "11", "100", "100", "111", '0', '-', "00"), -- i=10174
      ("1011111101000100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10175
      ("0101011101000000", '0', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10176
      ("0101111101000000", '1', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10177
      ("0101111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10178
      ("0100011101000000", '0', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10179
      ("0100111101000000", '1', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10180
      ("0100111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10181
      ("0000011111001000", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10182
      ("0000111111001000", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10183
      ("0000111111001000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10184
      ("1000011101000101", '0', '1', "00", "100", "101", "111", '0', '-', "00"), -- i=10185
      ("1000111101000101", '1', '1', "00", "100", "101", "111", '0', '-', "00"), -- i=10186
      ("1000111101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10187
      ("1001011101000101", '0', '1', "01", "100", "101", "111", '0', '-', "00"), -- i=10188
      ("1001111101000101", '1', '1', "01", "100", "101", "111", '0', '-', "00"), -- i=10189
      ("1001111101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10190
      ("1010011101000101", '0', '1', "10", "100", "101", "111", '0', '-', "00"), -- i=10191
      ("1010111101000101", '1', '1', "10", "100", "101", "111", '0', '-', "00"), -- i=10192
      ("1010111101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10193
      ("1011011101000101", '0', '1', "11", "100", "101", "111", '0', '-', "00"), -- i=10194
      ("1011111101000101", '1', '1', "11", "100", "101", "111", '0', '-', "00"), -- i=10195
      ("1011111101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10196
      ("0101011101000000", '0', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10197
      ("0101111101000000", '1', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10198
      ("0101111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10199
      ("0100011101000000", '0', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10200
      ("0100111101000000", '1', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10201
      ("0100111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10202
      ("0000011110001111", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10203
      ("0000111110001111", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10204
      ("0000111110001111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10205
      ("1000011101000110", '0', '1', "00", "100", "110", "111", '0', '-', "00"), -- i=10206
      ("1000111101000110", '1', '1', "00", "100", "110", "111", '0', '-', "00"), -- i=10207
      ("1000111101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10208
      ("1001011101000110", '0', '1', "01", "100", "110", "111", '0', '-', "00"), -- i=10209
      ("1001111101000110", '1', '1', "01", "100", "110", "111", '0', '-', "00"), -- i=10210
      ("1001111101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10211
      ("1010011101000110", '0', '1', "10", "100", "110", "111", '0', '-', "00"), -- i=10212
      ("1010111101000110", '1', '1', "10", "100", "110", "111", '0', '-', "00"), -- i=10213
      ("1010111101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10214
      ("1011011101000110", '0', '1', "11", "100", "110", "111", '0', '-', "00"), -- i=10215
      ("1011111101000110", '1', '1', "11", "100", "110", "111", '0', '-', "00"), -- i=10216
      ("1011111101000110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10217
      ("0101011101000000", '0', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10218
      ("0101111101000000", '1', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10219
      ("0101111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10220
      ("0100011101000000", '0', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10221
      ("0100111101000000", '1', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10222
      ("0100111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10223
      ("0000011101010010", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10224
      ("0000111101010010", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10225
      ("0000111101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10226
      ("1000011101000111", '0', '1', "00", "100", "111", "111", '0', '-', "00"), -- i=10227
      ("1000111101000111", '1', '1', "00", "100", "111", "111", '0', '-', "00"), -- i=10228
      ("1000111101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10229
      ("1001011101000111", '0', '1', "01", "100", "111", "111", '0', '-', "00"), -- i=10230
      ("1001111101000111", '1', '1', "01", "100", "111", "111", '0', '-', "00"), -- i=10231
      ("1001111101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10232
      ("1010011101000111", '0', '1', "10", "100", "111", "111", '0', '-', "00"), -- i=10233
      ("1010111101000111", '1', '1', "10", "100", "111", "111", '0', '-', "00"), -- i=10234
      ("1010111101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10235
      ("1011011101000111", '0', '1', "11", "100", "111", "111", '0', '-', "00"), -- i=10236
      ("1011111101000111", '1', '1', "11", "100", "111", "111", '0', '-', "00"), -- i=10237
      ("1011111101000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10238
      ("0101011101000000", '0', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10239
      ("0101111101000000", '1', '1', "--", "100", "---", "111", '0', '1', "01"), -- i=10240
      ("0101111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10241
      ("0100011101000000", '0', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10242
      ("0100111101000000", '1', '0', "--", "100", "111", "---", '1', '-', "--"), -- i=10243
      ("0100111101000000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10244
      ("0000011111101010", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10245
      ("0000111111101010", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10246
      ("0000111111101010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10247
      ("1000011101010000", '0', '1', "00", "101", "000", "111", '0', '-', "00"), -- i=10248
      ("1000111101010000", '1', '1', "00", "101", "000", "111", '0', '-', "00"), -- i=10249
      ("1000111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10250
      ("1001011101010000", '0', '1', "01", "101", "000", "111", '0', '-', "00"), -- i=10251
      ("1001111101010000", '1', '1', "01", "101", "000", "111", '0', '-', "00"), -- i=10252
      ("1001111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10253
      ("1010011101010000", '0', '1', "10", "101", "000", "111", '0', '-', "00"), -- i=10254
      ("1010111101010000", '1', '1', "10", "101", "000", "111", '0', '-', "00"), -- i=10255
      ("1010111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10256
      ("1011011101010000", '0', '1', "11", "101", "000", "111", '0', '-', "00"), -- i=10257
      ("1011111101010000", '1', '1', "11", "101", "000", "111", '0', '-', "00"), -- i=10258
      ("1011111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10259
      ("0101011101010000", '0', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10260
      ("0101111101010000", '1', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10261
      ("0101111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10262
      ("0100011101010000", '0', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10263
      ("0100111101010000", '1', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10264
      ("0100111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10265
      ("0000011110011111", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10266
      ("0000111110011111", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10267
      ("0000111110011111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10268
      ("1000011101010001", '0', '1', "00", "101", "001", "111", '0', '-', "00"), -- i=10269
      ("1000111101010001", '1', '1', "00", "101", "001", "111", '0', '-', "00"), -- i=10270
      ("1000111101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10271
      ("1001011101010001", '0', '1', "01", "101", "001", "111", '0', '-', "00"), -- i=10272
      ("1001111101010001", '1', '1', "01", "101", "001", "111", '0', '-', "00"), -- i=10273
      ("1001111101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10274
      ("1010011101010001", '0', '1', "10", "101", "001", "111", '0', '-', "00"), -- i=10275
      ("1010111101010001", '1', '1', "10", "101", "001", "111", '0', '-', "00"), -- i=10276
      ("1010111101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10277
      ("1011011101010001", '0', '1', "11", "101", "001", "111", '0', '-', "00"), -- i=10278
      ("1011111101010001", '1', '1', "11", "101", "001", "111", '0', '-', "00"), -- i=10279
      ("1011111101010001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10280
      ("0101011101010000", '0', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10281
      ("0101111101010000", '1', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10282
      ("0101111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10283
      ("0100011101010000", '0', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10284
      ("0100111101010000", '1', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10285
      ("0100111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10286
      ("0000011100111000", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10287
      ("0000111100111000", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10288
      ("0000111100111000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10289
      ("1000011101010010", '0', '1', "00", "101", "010", "111", '0', '-', "00"), -- i=10290
      ("1000111101010010", '1', '1', "00", "101", "010", "111", '0', '-', "00"), -- i=10291
      ("1000111101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10292
      ("1001011101010010", '0', '1', "01", "101", "010", "111", '0', '-', "00"), -- i=10293
      ("1001111101010010", '1', '1', "01", "101", "010", "111", '0', '-', "00"), -- i=10294
      ("1001111101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10295
      ("1010011101010010", '0', '1', "10", "101", "010", "111", '0', '-', "00"), -- i=10296
      ("1010111101010010", '1', '1', "10", "101", "010", "111", '0', '-', "00"), -- i=10297
      ("1010111101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10298
      ("1011011101010010", '0', '1', "11", "101", "010", "111", '0', '-', "00"), -- i=10299
      ("1011111101010010", '1', '1', "11", "101", "010", "111", '0', '-', "00"), -- i=10300
      ("1011111101010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10301
      ("0101011101010000", '0', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10302
      ("0101111101010000", '1', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10303
      ("0101111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10304
      ("0100011101010000", '0', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10305
      ("0100111101010000", '1', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10306
      ("0100111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10307
      ("0000011110110010", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10308
      ("0000111110110010", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10309
      ("0000111110110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10310
      ("1000011101010011", '0', '1', "00", "101", "011", "111", '0', '-', "00"), -- i=10311
      ("1000111101010011", '1', '1', "00", "101", "011", "111", '0', '-', "00"), -- i=10312
      ("1000111101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10313
      ("1001011101010011", '0', '1', "01", "101", "011", "111", '0', '-', "00"), -- i=10314
      ("1001111101010011", '1', '1', "01", "101", "011", "111", '0', '-', "00"), -- i=10315
      ("1001111101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10316
      ("1010011101010011", '0', '1', "10", "101", "011", "111", '0', '-', "00"), -- i=10317
      ("1010111101010011", '1', '1', "10", "101", "011", "111", '0', '-', "00"), -- i=10318
      ("1010111101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10319
      ("1011011101010011", '0', '1', "11", "101", "011", "111", '0', '-', "00"), -- i=10320
      ("1011111101010011", '1', '1', "11", "101", "011", "111", '0', '-', "00"), -- i=10321
      ("1011111101010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10322
      ("0101011101010000", '0', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10323
      ("0101111101010000", '1', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10324
      ("0101111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10325
      ("0100011101010000", '0', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10326
      ("0100111101010000", '1', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10327
      ("0100111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10328
      ("0000011111000111", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10329
      ("0000111111000111", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10330
      ("0000111111000111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10331
      ("1000011101010100", '0', '1', "00", "101", "100", "111", '0', '-', "00"), -- i=10332
      ("1000111101010100", '1', '1', "00", "101", "100", "111", '0', '-', "00"), -- i=10333
      ("1000111101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10334
      ("1001011101010100", '0', '1', "01", "101", "100", "111", '0', '-', "00"), -- i=10335
      ("1001111101010100", '1', '1', "01", "101", "100", "111", '0', '-', "00"), -- i=10336
      ("1001111101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10337
      ("1010011101010100", '0', '1', "10", "101", "100", "111", '0', '-', "00"), -- i=10338
      ("1010111101010100", '1', '1', "10", "101", "100", "111", '0', '-', "00"), -- i=10339
      ("1010111101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10340
      ("1011011101010100", '0', '1', "11", "101", "100", "111", '0', '-', "00"), -- i=10341
      ("1011111101010100", '1', '1', "11", "101", "100", "111", '0', '-', "00"), -- i=10342
      ("1011111101010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10343
      ("0101011101010000", '0', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10344
      ("0101111101010000", '1', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10345
      ("0101111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10346
      ("0100011101010000", '0', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10347
      ("0100111101010000", '1', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10348
      ("0100111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10349
      ("0000011101000101", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10350
      ("0000111101000101", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10351
      ("0000111101000101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10352
      ("1000011101010101", '0', '1', "00", "101", "101", "111", '0', '-', "00"), -- i=10353
      ("1000111101010101", '1', '1', "00", "101", "101", "111", '0', '-', "00"), -- i=10354
      ("1000111101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10355
      ("1001011101010101", '0', '1', "01", "101", "101", "111", '0', '-', "00"), -- i=10356
      ("1001111101010101", '1', '1', "01", "101", "101", "111", '0', '-', "00"), -- i=10357
      ("1001111101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10358
      ("1010011101010101", '0', '1', "10", "101", "101", "111", '0', '-', "00"), -- i=10359
      ("1010111101010101", '1', '1', "10", "101", "101", "111", '0', '-', "00"), -- i=10360
      ("1010111101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10361
      ("1011011101010101", '0', '1', "11", "101", "101", "111", '0', '-', "00"), -- i=10362
      ("1011111101010101", '1', '1', "11", "101", "101", "111", '0', '-', "00"), -- i=10363
      ("1011111101010101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10364
      ("0101011101010000", '0', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10365
      ("0101111101010000", '1', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10366
      ("0101111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10367
      ("0100011101010000", '0', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10368
      ("0100111101010000", '1', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10369
      ("0100111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10370
      ("0000011111010010", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10371
      ("0000111111010010", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10372
      ("0000111111010010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10373
      ("1000011101010110", '0', '1', "00", "101", "110", "111", '0', '-', "00"), -- i=10374
      ("1000111101010110", '1', '1', "00", "101", "110", "111", '0', '-', "00"), -- i=10375
      ("1000111101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10376
      ("1001011101010110", '0', '1', "01", "101", "110", "111", '0', '-', "00"), -- i=10377
      ("1001111101010110", '1', '1', "01", "101", "110", "111", '0', '-', "00"), -- i=10378
      ("1001111101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10379
      ("1010011101010110", '0', '1', "10", "101", "110", "111", '0', '-', "00"), -- i=10380
      ("1010111101010110", '1', '1', "10", "101", "110", "111", '0', '-', "00"), -- i=10381
      ("1010111101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10382
      ("1011011101010110", '0', '1', "11", "101", "110", "111", '0', '-', "00"), -- i=10383
      ("1011111101010110", '1', '1', "11", "101", "110", "111", '0', '-', "00"), -- i=10384
      ("1011111101010110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10385
      ("0101011101010000", '0', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10386
      ("0101111101010000", '1', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10387
      ("0101111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10388
      ("0100011101010000", '0', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10389
      ("0100111101010000", '1', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10390
      ("0100111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10391
      ("0000011111011010", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10392
      ("0000111111011010", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10393
      ("0000111111011010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10394
      ("1000011101010111", '0', '1', "00", "101", "111", "111", '0', '-', "00"), -- i=10395
      ("1000111101010111", '1', '1', "00", "101", "111", "111", '0', '-', "00"), -- i=10396
      ("1000111101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10397
      ("1001011101010111", '0', '1', "01", "101", "111", "111", '0', '-', "00"), -- i=10398
      ("1001111101010111", '1', '1', "01", "101", "111", "111", '0', '-', "00"), -- i=10399
      ("1001111101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10400
      ("1010011101010111", '0', '1', "10", "101", "111", "111", '0', '-', "00"), -- i=10401
      ("1010111101010111", '1', '1', "10", "101", "111", "111", '0', '-', "00"), -- i=10402
      ("1010111101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10403
      ("1011011101010111", '0', '1', "11", "101", "111", "111", '0', '-', "00"), -- i=10404
      ("1011111101010111", '1', '1', "11", "101", "111", "111", '0', '-', "00"), -- i=10405
      ("1011111101010111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10406
      ("0101011101010000", '0', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10407
      ("0101111101010000", '1', '1', "--", "101", "---", "111", '0', '1', "01"), -- i=10408
      ("0101111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10409
      ("0100011101010000", '0', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10410
      ("0100111101010000", '1', '0', "--", "101", "111", "---", '1', '-', "--"), -- i=10411
      ("0100111101010000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10412
      ("0000011110110111", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10413
      ("0000111110110111", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10414
      ("0000111110110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10415
      ("1000011101100000", '0', '1', "00", "110", "000", "111", '0', '-', "00"), -- i=10416
      ("1000111101100000", '1', '1', "00", "110", "000", "111", '0', '-', "00"), -- i=10417
      ("1000111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10418
      ("1001011101100000", '0', '1', "01", "110", "000", "111", '0', '-', "00"), -- i=10419
      ("1001111101100000", '1', '1', "01", "110", "000", "111", '0', '-', "00"), -- i=10420
      ("1001111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10421
      ("1010011101100000", '0', '1', "10", "110", "000", "111", '0', '-', "00"), -- i=10422
      ("1010111101100000", '1', '1', "10", "110", "000", "111", '0', '-', "00"), -- i=10423
      ("1010111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10424
      ("1011011101100000", '0', '1', "11", "110", "000", "111", '0', '-', "00"), -- i=10425
      ("1011111101100000", '1', '1', "11", "110", "000", "111", '0', '-', "00"), -- i=10426
      ("1011111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10427
      ("0101011101100000", '0', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10428
      ("0101111101100000", '1', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10429
      ("0101111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10430
      ("0100011101100000", '0', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10431
      ("0100111101100000", '1', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10432
      ("0100111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10433
      ("0000011111010100", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10434
      ("0000111111010100", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10435
      ("0000111111010100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10436
      ("1000011101100001", '0', '1', "00", "110", "001", "111", '0', '-', "00"), -- i=10437
      ("1000111101100001", '1', '1', "00", "110", "001", "111", '0', '-', "00"), -- i=10438
      ("1000111101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10439
      ("1001011101100001", '0', '1', "01", "110", "001", "111", '0', '-', "00"), -- i=10440
      ("1001111101100001", '1', '1', "01", "110", "001", "111", '0', '-', "00"), -- i=10441
      ("1001111101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10442
      ("1010011101100001", '0', '1', "10", "110", "001", "111", '0', '-', "00"), -- i=10443
      ("1010111101100001", '1', '1', "10", "110", "001", "111", '0', '-', "00"), -- i=10444
      ("1010111101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10445
      ("1011011101100001", '0', '1', "11", "110", "001", "111", '0', '-', "00"), -- i=10446
      ("1011111101100001", '1', '1', "11", "110", "001", "111", '0', '-', "00"), -- i=10447
      ("1011111101100001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10448
      ("0101011101100000", '0', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10449
      ("0101111101100000", '1', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10450
      ("0101111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10451
      ("0100011101100000", '0', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10452
      ("0100111101100000", '1', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10453
      ("0100111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10454
      ("0000011100010011", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10455
      ("0000111100010011", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10456
      ("0000111100010011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10457
      ("1000011101100010", '0', '1', "00", "110", "010", "111", '0', '-', "00"), -- i=10458
      ("1000111101100010", '1', '1', "00", "110", "010", "111", '0', '-', "00"), -- i=10459
      ("1000111101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10460
      ("1001011101100010", '0', '1', "01", "110", "010", "111", '0', '-', "00"), -- i=10461
      ("1001111101100010", '1', '1', "01", "110", "010", "111", '0', '-', "00"), -- i=10462
      ("1001111101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10463
      ("1010011101100010", '0', '1', "10", "110", "010", "111", '0', '-', "00"), -- i=10464
      ("1010111101100010", '1', '1', "10", "110", "010", "111", '0', '-', "00"), -- i=10465
      ("1010111101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10466
      ("1011011101100010", '0', '1', "11", "110", "010", "111", '0', '-', "00"), -- i=10467
      ("1011111101100010", '1', '1', "11", "110", "010", "111", '0', '-', "00"), -- i=10468
      ("1011111101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10469
      ("0101011101100000", '0', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10470
      ("0101111101100000", '1', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10471
      ("0101111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10472
      ("0100011101100000", '0', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10473
      ("0100111101100000", '1', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10474
      ("0100111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10475
      ("0000011101111110", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10476
      ("0000111101111110", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10477
      ("0000111101111110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10478
      ("1000011101100011", '0', '1', "00", "110", "011", "111", '0', '-', "00"), -- i=10479
      ("1000111101100011", '1', '1', "00", "110", "011", "111", '0', '-', "00"), -- i=10480
      ("1000111101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10481
      ("1001011101100011", '0', '1', "01", "110", "011", "111", '0', '-', "00"), -- i=10482
      ("1001111101100011", '1', '1', "01", "110", "011", "111", '0', '-', "00"), -- i=10483
      ("1001111101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10484
      ("1010011101100011", '0', '1', "10", "110", "011", "111", '0', '-', "00"), -- i=10485
      ("1010111101100011", '1', '1', "10", "110", "011", "111", '0', '-', "00"), -- i=10486
      ("1010111101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10487
      ("1011011101100011", '0', '1', "11", "110", "011", "111", '0', '-', "00"), -- i=10488
      ("1011111101100011", '1', '1', "11", "110", "011", "111", '0', '-', "00"), -- i=10489
      ("1011111101100011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10490
      ("0101011101100000", '0', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10491
      ("0101111101100000", '1', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10492
      ("0101111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10493
      ("0100011101100000", '0', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10494
      ("0100111101100000", '1', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10495
      ("0100111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10496
      ("0000011101110111", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10497
      ("0000111101110111", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10498
      ("0000111101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10499
      ("1000011101100100", '0', '1', "00", "110", "100", "111", '0', '-', "00"), -- i=10500
      ("1000111101100100", '1', '1', "00", "110", "100", "111", '0', '-', "00"), -- i=10501
      ("1000111101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10502
      ("1001011101100100", '0', '1', "01", "110", "100", "111", '0', '-', "00"), -- i=10503
      ("1001111101100100", '1', '1', "01", "110", "100", "111", '0', '-', "00"), -- i=10504
      ("1001111101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10505
      ("1010011101100100", '0', '1', "10", "110", "100", "111", '0', '-', "00"), -- i=10506
      ("1010111101100100", '1', '1', "10", "110", "100", "111", '0', '-', "00"), -- i=10507
      ("1010111101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10508
      ("1011011101100100", '0', '1', "11", "110", "100", "111", '0', '-', "00"), -- i=10509
      ("1011111101100100", '1', '1', "11", "110", "100", "111", '0', '-', "00"), -- i=10510
      ("1011111101100100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10511
      ("0101011101100000", '0', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10512
      ("0101111101100000", '1', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10513
      ("0101111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10514
      ("0100011101100000", '0', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10515
      ("0100111101100000", '1', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10516
      ("0100111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10517
      ("0000011101001100", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10518
      ("0000111101001100", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10519
      ("0000111101001100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10520
      ("1000011101100101", '0', '1', "00", "110", "101", "111", '0', '-', "00"), -- i=10521
      ("1000111101100101", '1', '1', "00", "110", "101", "111", '0', '-', "00"), -- i=10522
      ("1000111101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10523
      ("1001011101100101", '0', '1', "01", "110", "101", "111", '0', '-', "00"), -- i=10524
      ("1001111101100101", '1', '1', "01", "110", "101", "111", '0', '-', "00"), -- i=10525
      ("1001111101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10526
      ("1010011101100101", '0', '1', "10", "110", "101", "111", '0', '-', "00"), -- i=10527
      ("1010111101100101", '1', '1', "10", "110", "101", "111", '0', '-', "00"), -- i=10528
      ("1010111101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10529
      ("1011011101100101", '0', '1', "11", "110", "101", "111", '0', '-', "00"), -- i=10530
      ("1011111101100101", '1', '1', "11", "110", "101", "111", '0', '-', "00"), -- i=10531
      ("1011111101100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10532
      ("0101011101100000", '0', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10533
      ("0101111101100000", '1', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10534
      ("0101111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10535
      ("0100011101100000", '0', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10536
      ("0100111101100000", '1', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10537
      ("0100111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10538
      ("0000011101011011", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10539
      ("0000111101011011", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10540
      ("0000111101011011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10541
      ("1000011101100110", '0', '1', "00", "110", "110", "111", '0', '-', "00"), -- i=10542
      ("1000111101100110", '1', '1', "00", "110", "110", "111", '0', '-', "00"), -- i=10543
      ("1000111101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10544
      ("1001011101100110", '0', '1', "01", "110", "110", "111", '0', '-', "00"), -- i=10545
      ("1001111101100110", '1', '1', "01", "110", "110", "111", '0', '-', "00"), -- i=10546
      ("1001111101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10547
      ("1010011101100110", '0', '1', "10", "110", "110", "111", '0', '-', "00"), -- i=10548
      ("1010111101100110", '1', '1', "10", "110", "110", "111", '0', '-', "00"), -- i=10549
      ("1010111101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10550
      ("1011011101100110", '0', '1', "11", "110", "110", "111", '0', '-', "00"), -- i=10551
      ("1011111101100110", '1', '1', "11", "110", "110", "111", '0', '-', "00"), -- i=10552
      ("1011111101100110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10553
      ("0101011101100000", '0', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10554
      ("0101111101100000", '1', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10555
      ("0101111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10556
      ("0100011101100000", '0', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10557
      ("0100111101100000", '1', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10558
      ("0100111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10559
      ("0000011110100101", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10560
      ("0000111110100101", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10561
      ("0000111110100101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10562
      ("1000011101100111", '0', '1', "00", "110", "111", "111", '0', '-', "00"), -- i=10563
      ("1000111101100111", '1', '1', "00", "110", "111", "111", '0', '-', "00"), -- i=10564
      ("1000111101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10565
      ("1001011101100111", '0', '1', "01", "110", "111", "111", '0', '-', "00"), -- i=10566
      ("1001111101100111", '1', '1', "01", "110", "111", "111", '0', '-', "00"), -- i=10567
      ("1001111101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10568
      ("1010011101100111", '0', '1', "10", "110", "111", "111", '0', '-', "00"), -- i=10569
      ("1010111101100111", '1', '1', "10", "110", "111", "111", '0', '-', "00"), -- i=10570
      ("1010111101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10571
      ("1011011101100111", '0', '1', "11", "110", "111", "111", '0', '-', "00"), -- i=10572
      ("1011111101100111", '1', '1', "11", "110", "111", "111", '0', '-', "00"), -- i=10573
      ("1011111101100111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10574
      ("0101011101100000", '0', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10575
      ("0101111101100000", '1', '1', "--", "110", "---", "111", '0', '1', "01"), -- i=10576
      ("0101111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10577
      ("0100011101100000", '0', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10578
      ("0100111101100000", '1', '0', "--", "110", "111", "---", '1', '-', "--"), -- i=10579
      ("0100111101100000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10580
      ("0000011110001100", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10581
      ("0000111110001100", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10582
      ("0000111110001100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10583
      ("1000011101110000", '0', '1', "00", "111", "000", "111", '0', '-', "00"), -- i=10584
      ("1000111101110000", '1', '1', "00", "111", "000", "111", '0', '-', "00"), -- i=10585
      ("1000111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10586
      ("1001011101110000", '0', '1', "01", "111", "000", "111", '0', '-', "00"), -- i=10587
      ("1001111101110000", '1', '1', "01", "111", "000", "111", '0', '-', "00"), -- i=10588
      ("1001111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10589
      ("1010011101110000", '0', '1', "10", "111", "000", "111", '0', '-', "00"), -- i=10590
      ("1010111101110000", '1', '1', "10", "111", "000", "111", '0', '-', "00"), -- i=10591
      ("1010111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10592
      ("1011011101110000", '0', '1', "11", "111", "000", "111", '0', '-', "00"), -- i=10593
      ("1011111101110000", '1', '1', "11", "111", "000", "111", '0', '-', "00"), -- i=10594
      ("1011111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10595
      ("0101011101110000", '0', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10596
      ("0101111101110000", '1', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10597
      ("0101111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10598
      ("0100011101110000", '0', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10599
      ("0100111101110000", '1', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10600
      ("0100111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10601
      ("0000011100111011", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10602
      ("0000111100111011", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10603
      ("0000111100111011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10604
      ("1000011101110001", '0', '1', "00", "111", "001", "111", '0', '-', "00"), -- i=10605
      ("1000111101110001", '1', '1', "00", "111", "001", "111", '0', '-', "00"), -- i=10606
      ("1000111101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10607
      ("1001011101110001", '0', '1', "01", "111", "001", "111", '0', '-', "00"), -- i=10608
      ("1001111101110001", '1', '1', "01", "111", "001", "111", '0', '-', "00"), -- i=10609
      ("1001111101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10610
      ("1010011101110001", '0', '1', "10", "111", "001", "111", '0', '-', "00"), -- i=10611
      ("1010111101110001", '1', '1', "10", "111", "001", "111", '0', '-', "00"), -- i=10612
      ("1010111101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10613
      ("1011011101110001", '0', '1', "11", "111", "001", "111", '0', '-', "00"), -- i=10614
      ("1011111101110001", '1', '1', "11", "111", "001", "111", '0', '-', "00"), -- i=10615
      ("1011111101110001", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10616
      ("0101011101110000", '0', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10617
      ("0101111101110000", '1', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10618
      ("0101111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10619
      ("0100011101110000", '0', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10620
      ("0100111101110000", '1', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10621
      ("0100111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10622
      ("0000011101001000", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10623
      ("0000111101001000", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10624
      ("0000111101001000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10625
      ("1000011101110010", '0', '1', "00", "111", "010", "111", '0', '-', "00"), -- i=10626
      ("1000111101110010", '1', '1', "00", "111", "010", "111", '0', '-', "00"), -- i=10627
      ("1000111101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10628
      ("1001011101110010", '0', '1', "01", "111", "010", "111", '0', '-', "00"), -- i=10629
      ("1001111101110010", '1', '1', "01", "111", "010", "111", '0', '-', "00"), -- i=10630
      ("1001111101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10631
      ("1010011101110010", '0', '1', "10", "111", "010", "111", '0', '-', "00"), -- i=10632
      ("1010111101110010", '1', '1', "10", "111", "010", "111", '0', '-', "00"), -- i=10633
      ("1010111101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10634
      ("1011011101110010", '0', '1', "11", "111", "010", "111", '0', '-', "00"), -- i=10635
      ("1011111101110010", '1', '1', "11", "111", "010", "111", '0', '-', "00"), -- i=10636
      ("1011111101110010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10637
      ("0101011101110000", '0', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10638
      ("0101111101110000", '1', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10639
      ("0101111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10640
      ("0100011101110000", '0', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10641
      ("0100111101110000", '1', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10642
      ("0100111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10643
      ("0000011111011000", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10644
      ("0000111111011000", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10645
      ("0000111111011000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10646
      ("1000011101110011", '0', '1', "00", "111", "011", "111", '0', '-', "00"), -- i=10647
      ("1000111101110011", '1', '1', "00", "111", "011", "111", '0', '-', "00"), -- i=10648
      ("1000111101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10649
      ("1001011101110011", '0', '1', "01", "111", "011", "111", '0', '-', "00"), -- i=10650
      ("1001111101110011", '1', '1', "01", "111", "011", "111", '0', '-', "00"), -- i=10651
      ("1001111101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10652
      ("1010011101110011", '0', '1', "10", "111", "011", "111", '0', '-', "00"), -- i=10653
      ("1010111101110011", '1', '1', "10", "111", "011", "111", '0', '-', "00"), -- i=10654
      ("1010111101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10655
      ("1011011101110011", '0', '1', "11", "111", "011", "111", '0', '-', "00"), -- i=10656
      ("1011111101110011", '1', '1', "11", "111", "011", "111", '0', '-', "00"), -- i=10657
      ("1011111101110011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10658
      ("0101011101110000", '0', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10659
      ("0101111101110000", '1', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10660
      ("0101111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10661
      ("0100011101110000", '0', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10662
      ("0100111101110000", '1', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10663
      ("0100111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10664
      ("0000011100011101", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10665
      ("0000111100011101", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10666
      ("0000111100011101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10667
      ("1000011101110100", '0', '1', "00", "111", "100", "111", '0', '-', "00"), -- i=10668
      ("1000111101110100", '1', '1', "00", "111", "100", "111", '0', '-', "00"), -- i=10669
      ("1000111101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10670
      ("1001011101110100", '0', '1', "01", "111", "100", "111", '0', '-', "00"), -- i=10671
      ("1001111101110100", '1', '1', "01", "111", "100", "111", '0', '-', "00"), -- i=10672
      ("1001111101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10673
      ("1010011101110100", '0', '1', "10", "111", "100", "111", '0', '-', "00"), -- i=10674
      ("1010111101110100", '1', '1', "10", "111", "100", "111", '0', '-', "00"), -- i=10675
      ("1010111101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10676
      ("1011011101110100", '0', '1', "11", "111", "100", "111", '0', '-', "00"), -- i=10677
      ("1011111101110100", '1', '1', "11", "111", "100", "111", '0', '-', "00"), -- i=10678
      ("1011111101110100", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10679
      ("0101011101110000", '0', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10680
      ("0101111101110000", '1', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10681
      ("0101111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10682
      ("0100011101110000", '0', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10683
      ("0100111101110000", '1', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10684
      ("0100111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10685
      ("0000011101011010", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10686
      ("0000111101011010", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10687
      ("0000111101011010", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10688
      ("1000011101110101", '0', '1', "00", "111", "101", "111", '0', '-', "00"), -- i=10689
      ("1000111101110101", '1', '1', "00", "111", "101", "111", '0', '-', "00"), -- i=10690
      ("1000111101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10691
      ("1001011101110101", '0', '1', "01", "111", "101", "111", '0', '-', "00"), -- i=10692
      ("1001111101110101", '1', '1', "01", "111", "101", "111", '0', '-', "00"), -- i=10693
      ("1001111101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10694
      ("1010011101110101", '0', '1', "10", "111", "101", "111", '0', '-', "00"), -- i=10695
      ("1010111101110101", '1', '1', "10", "111", "101", "111", '0', '-', "00"), -- i=10696
      ("1010111101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10697
      ("1011011101110101", '0', '1', "11", "111", "101", "111", '0', '-', "00"), -- i=10698
      ("1011111101110101", '1', '1', "11", "111", "101", "111", '0', '-', "00"), -- i=10699
      ("1011111101110101", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10700
      ("0101011101110000", '0', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10701
      ("0101111101110000", '1', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10702
      ("0101111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10703
      ("0100011101110000", '0', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10704
      ("0100111101110000", '1', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10705
      ("0100111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10706
      ("0000011100001110", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10707
      ("0000111100001110", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10708
      ("0000111100001110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10709
      ("1000011101110110", '0', '1', "00", "111", "110", "111", '0', '-', "00"), -- i=10710
      ("1000111101110110", '1', '1', "00", "111", "110", "111", '0', '-', "00"), -- i=10711
      ("1000111101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10712
      ("1001011101110110", '0', '1', "01", "111", "110", "111", '0', '-', "00"), -- i=10713
      ("1001111101110110", '1', '1', "01", "111", "110", "111", '0', '-', "00"), -- i=10714
      ("1001111101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10715
      ("1010011101110110", '0', '1', "10", "111", "110", "111", '0', '-', "00"), -- i=10716
      ("1010111101110110", '1', '1', "10", "111", "110", "111", '0', '-', "00"), -- i=10717
      ("1010111101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10718
      ("1011011101110110", '0', '1', "11", "111", "110", "111", '0', '-', "00"), -- i=10719
      ("1011111101110110", '1', '1', "11", "111", "110", "111", '0', '-', "00"), -- i=10720
      ("1011111101110110", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10721
      ("0101011101110000", '0', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10722
      ("0101111101110000", '1', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10723
      ("0101111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10724
      ("0100011101110000", '0', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10725
      ("0100111101110000", '1', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10726
      ("0100111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10727
      ("0000011101000011", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10728
      ("0000111101000011", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10729
      ("0000111101000011", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10730
      ("1000011101110111", '0', '1', "00", "111", "111", "111", '0', '-', "00"), -- i=10731
      ("1000111101110111", '1', '1', "00", "111", "111", "111", '0', '-', "00"), -- i=10732
      ("1000111101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10733
      ("1001011101110111", '0', '1', "01", "111", "111", "111", '0', '-', "00"), -- i=10734
      ("1001111101110111", '1', '1', "01", "111", "111", "111", '0', '-', "00"), -- i=10735
      ("1001111101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10736
      ("1010011101110111", '0', '1', "10", "111", "111", "111", '0', '-', "00"), -- i=10737
      ("1010111101110111", '1', '1', "10", "111", "111", "111", '0', '-', "00"), -- i=10738
      ("1010111101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10739
      ("1011011101110111", '0', '1', "11", "111", "111", "111", '0', '-', "00"), -- i=10740
      ("1011111101110111", '1', '1', "11", "111", "111", "111", '0', '-', "00"), -- i=10741
      ("1011111101110111", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10742
      ("0101011101110000", '0', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10743
      ("0101111101110000", '1', '1', "--", "111", "---", "111", '0', '1', "01"), -- i=10744
      ("0101111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10745
      ("0100011101110000", '0', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10746
      ("0100111101110000", '1', '0', "--", "111", "111", "---", '1', '-', "--"), -- i=10747
      ("0100111101110000", '0', '0', "00", "000", "000", "000", '0', '0', "00"), -- i=10748
      ("0000011101100010", '0', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10749
      ("0000111101100010", '1', '1', "--", "---", "---", "111", '0', '-', "10"), -- i=10750
      ("0000111101100010", '0', '0', "00", "000", "000", "000", '0', '0', "00"));
  begin
    for i in patterns'range loop
      INST <= patterns(i).INST;
      FL_Z <= patterns(i).FL_Z;
      wait for 10 ns;
      assert std_match(ALUOP, patterns(i).ALUOP) OR (ALUOP = "ZZ" AND patterns(i).ALUOP = "ZZ")
        report "wrong value for ALUOP, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).ALUOP) & ", found " & to_string(ALUOP) severity error;assert std_match(RS1, patterns(i).RS1) OR (RS1 = "ZZZ" AND patterns(i).RS1 = "ZZZ")
        report "wrong value for RS1, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).RS1) & ", found " & to_string(RS1) severity error;assert std_match(RS2, patterns(i).RS2) OR (RS2 = "ZZZ" AND patterns(i).RS2 = "ZZZ")
        report "wrong value for RS2, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).RS2) & ", found " & to_string(RS2) severity error;assert std_match(WS, patterns(i).WS) OR (WS = "ZZZ" AND patterns(i).WS = "ZZZ")
        report "wrong value for WS, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).WS) & ", found " & to_string(WS) severity error;assert std_match(STR, patterns(i).STR) OR (STR = 'Z' AND patterns(i).STR = 'Z')
        report "wrong value for STR, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).STR) & ", found " & std_logic'image(STR) severity error;assert std_match(WE, patterns(i).WE) OR (WE = 'Z' AND patterns(i).WE = 'Z')
        report "wrong value for WE, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).WE) & ", found " & std_logic'image(WE) severity error;assert std_match(DMUX, patterns(i).DMUX) OR (DMUX = "ZZ" AND patterns(i).DMUX = "ZZ")
        report "wrong value for DMUX, i=" & integer'image(i)
         & ", expected " & to_string(patterns(i).DMUX) & ", found " & to_string(DMUX) severity error;assert std_match(LDR, patterns(i).LDR) OR (LDR = 'Z' AND patterns(i).LDR = 'Z')
        report "wrong value for LDR, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).LDR) & ", found " & std_logic'image(LDR) severity error;assert std_match(FL_EN, patterns(i).FL_EN) OR (FL_EN = 'Z' AND patterns(i).FL_EN = 'Z')
        report "wrong value for FL_EN, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).FL_EN) & ", found " & std_logic'image(FL_EN) severity error;assert std_match(HE, patterns(i).HE) OR (HE = 'Z' AND patterns(i).HE = 'Z')
        report "wrong value for HE, i=" & integer'image(i)
         & ", expected " & std_logic'image(patterns(i).HE) & ", found " & std_logic'image(HE) severity error;end loop;
    wait;
  end process;
end behav;
